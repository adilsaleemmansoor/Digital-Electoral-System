PK   ���X�v�[E7  `�    cirkitFile.json�}���6��(��v�w�c|;�]����j�v��t�IR*>�XY:Wұ��A�3�M�ґ���������m��������&���6}/֋|���b�[n�WY0�z�n�������f�^�7����۫���;��7�ɶ"-���(��䂅��!w|^DN���i�e9K�<_�����ϧ#0cw��9�"�n���]x�L܅o���]�L�Eh���]D�L�El���]$�L��2w����U��Jf�,�!$swi!Y�;Lc���eCH�N�B�0w������4��,�]�1��[��Nc���wCH��������B�0�������4��,�}�1�da�;�!$s�i!Y���!�T��_��D�t|��N�e�x�W�Y\�%��I��9�À�#r0E�ωL�s"S�:>?��7�n6k��/x���ㆾ+-2I��K3GE즮(���2�y����u��rE٬��r��Y����	�tL�D��i"S��4��)�`�����]W1���34|>��@��|B�rTB�C�P����|��5PY�C�*S��t����rӟ���YM�����#��i*�d(�Aea>��<�s^���P΃�0����}�P΃��܇�<�,�}�P΃��܇�<�,�g�C9*s�9��0���9������H-k8�7�N��fp��n�,Ŀ�1�/l2����s�w�a�X�]�NiT�I�s'����K�;�w��2?E�nx�Z6��gx�8��q���cXv���j�a�k��1���'n�D<b�Ɖ��^�0�SOd�<�k_�d&fϝ{��D�1{Ǡ�ZyZӋ��X������څX��������EX���������X�����H��%X����{��c7,����ER�H
ʏ����E`��q��S����c,?��Ё�GX~�O�[��6����{�V�8���k�E5�^p���Q��So����#,?��]��GX~�O�u������S�`�����S�`���U�/V���`�10?U]�`�10?U�`�10?U��`�10?U��`�10?UE���u��K��k�͸A�8�i^��h��*O���E�8Y�%��GNR��#������_��ҷ.m2�ޚ�'�ě�gX��"�+�ۃ�Z#�j�;5���c����ײ��!����ײQ?��jG�g���b����W���!����*;�M��L*j��Pʎ^�F���5�~Q��ʎ^����ʎ^�F���5Z�~���ʎ^����ʎ^�F��<����5j�&�`6R��ؖ�� X~th��m���dlD?p|��Q�6�8����(i����`�i��M����V��4J�&�A�G,m~F�wh:|�Cr�y���ਇ\q6�8���Ө�����`�iT�M��d�����FE�<�~���O�"nD?��p�B�8����`�iT�M���_��4*�&�A��/X~q� ���,?���	x�����FE�<�~���O��mD?p�1T�f^�x��T�Ux%O��ee&��{~�xY�eXE�^	_�{sK����'5�7׍<uyX��NY:>�����<�B��h��I����Խ��I���=��� vr���^�:	�K'c���Ћ<��vR��k'u�vR��k'֕>~	��#QaW&�-'&��F��MN�o@�B[s�?���orj�{��Ss��( q�E�~K��$i.�+��藮��~*��XD�W��G�������!�w�8@�n���� �{�8@\(���\�S@\(Ƥ�) 1i.��ٽ�b�f��R˚ݛk$����`�4�v���o�<�����#�ɩ�S3�S�|�Ã��c�������ֶ��M����0i%]#�ɩ��;����-&��|�l�fr�����L���������N�MN������<C����$t˔��a\��x*y#|9YE�恗�C9R���ga�KI7I3��c�K�	3'�� 2V�I:tvJ���g��G<w^��$�N�
5X��[!� 8;�{�ى>�$��z��82����Q#.�nUx��q�{��H�Ĥ���S���,��j��z�K�+�n�r���On���dNk\P�9-��ڪ�Tm\�a����0U��b����e1�@@�N�F �j�Y#P�-��ޓ�"q^�a~��7
��5�	��y���eA�`���8
����	��̉���`A�`~���8
���	7��M�a~���8
��G�	��9̏���=fA�`~���8
���	��9̏���0@�
5��b��P�Ũ(F�n����Q�tV�yfƨbq�ŗ��q�K]�
�Ѹå��b4�n�k+��;[�E(F WKɡ�߀VH,����c�2�g`:�7
��C!/��4>c&/6�s�(�c�,/��B�ss�($R����̍��H9�*0N0?�B"�P�_��8��8
��C!u���($R��u0�̏��H9�W�0N0?އ�[$��c �Z}��@m�p���O�����ͥ`0�6�����е��ks���ͅb0�����t �@s�8*P�6W����"쵹�F���2]mpmoV�Q�������0
4����u����MF���4pT��6���0�(�\��
������K��Q������� 4��p�6 E6�vl� �R�e)���c��v�� �^V�vl���Ejk�m�^	 �`��	@"�	�����N���Nf�m�VxX��vB1+l;�Q��"���Ya۱������
ێ��Hm�eV�v�̀�E�Y��Ya۱o�����
ێ=�Hm-�����S��"���Ya۱�����
ێ}"�Hm��eV�v�!��Ejk'.�¶c	<,R[;q��{O�a�ڶ�"J<���ؗ�Զ��m��`���Z�i���
��U�hε�>��f���
��U�F���u��U�>��հ]5c��Vt��U�>Q���]���qK3��G�j��v}"�;t+�j�3�Oݭ�j��v}�>*PW\���kX�U3��.;`EW\���Q����]�H^��N``#�ѯO� ��V�M�Ejk)�w�V�M�Ejk'���V�>q,R[;�����`���	���կO� ���Nf��~}�X��vB���y��`L�⏼��m��c�`���	ɬ�կO� ���NXf��~}�X�;q�����`��ډˬ�կO� ����+1;q�n��X��v�2+l��'�"���Ya�_�8�����
[���	�Hm��eV���'N�Ejk'.��V�>q,R[;q�����`��ډ�:ض�O��^�!a���$j�:����iP�eQD��Fh���5��ҳ:�&J�z�'���eθ�j8�	�I|�sDz�W�nDх�2�	eTʨ.A�����L�xa�$�/���"
B/�b\ʨ.$�Q]H(���6�vǞF�6�%	\�KP����xݹ�JyR��IrWm[�|'+�l�{A�Ǣ(��%���^�놑
�G$�Q]�<�E�ikRS�t}'�S��ce^�n-zv~�D�t)K�������3MB}�i;CPF�i�?f/$�`�N�PzV��D�Y�Z�g5iM����u�d���ۨDc��v CΗ�y_Ƅ�}2�����-ta0Vܷ��.��a�3���89�{f342�����HӅ9Xqs�']�����^6�0��T����;i�.Ɗ�Q+NB�Ly)ƅ�s#OE>2�I�P�nxII�TH(�\�0㥼�$�|ǏY.��0s2/�@Fy��PPF�d��G<w^�����u�T��l꺅��q.$�Q."-O�ԉx�?�e��z��d��,�G3�!ABac����76g$�����Y�7��>݋����`�7AU����~������
�7�0��B���G!�@@���F �z�Q#P��(���p�To8
a�7�06ŸH��ƹm��f0ǍB:l8�����QH�G1�`���8
��(�̇3�G!6�p��q��(�Æ�N��7n����QH�G1�`~���8
��(�̏s�G!6�p��q��$��[ J��}	���C�=���]�*F(F�N����Ѹ˥���b4�p�kΠ��[�j-(F�Ζ��	���Rr(��;`.�qn�	��J0N0׍B"�P�+�8��7
��C!��s�($R��e4�̍��H9�0N0?�B"�P�_~�8��8
��C!i���($R��e�̏��H9�T0N0?އ��2|ku4j�� �cQt4*�kǢ�hT��6�v,�Q��������Ch���F�j�kǢ�Z�)�Q����ڱ(:D��J
hT��6�v,�Q��������Ch���F�j�kǢ�Z�'�Q����ڱ(:D���	hT��6�v,�����	��ˌc��vB.+l�E��"��vى��ˌ�a���	����Z���N�e�mע�pX��vB0+l�E��"���Ya۵(:���P�
ۮE��Hm�cV�v-��Ejk'$�¶kQt8,R[;a��]���a�o��eV�v-��Ejk'.�¶kQt8,R[K����e�e��Hm��eV�v-��Ejk'.�¶kQt8,R[;q��]���a��ډˬ��Z���N\f�mע�pX��v�2+l�E��"���鲥~�GV�U�>Q��f���
��W��Dj��]5�j�]mpծO�G�j��v}"��g+�j�5�ϫ��j��v}�>*PW\���ߡ[�U3��~�nEW\���Q����]�H]����qu�+���]���
��W��D��v;������u&�hk)�vى�t+�&�"��zYa�_�8�����
[���	�Hm�`V���'N�Ejk'��V�>q,R[;������`���	Ǭ�կO� ���NHf��~}�X��v�2+l��'�"�,؉ˬ�կO� ���N\f��~}�X���^�ى�t+�&�"���Ya�_�8�����
[���	�Hm��eV���'N�Ejk'.��V�>q,R[;q�����`��ډˬ�կO� ���N\Fb{���J�	ee&Q�ԉ=�p��H�2,�"��7B�g�YM���a5Qz�s=��<,s���q��L�N⻞#���"t#�.$�Q]H(���PFu	���,���g�S'�~�d�Qz��㺐PFu!���BB�%b�_a�d�%���(#G$q�Q�?�	eTʨ.$�Q]Ҩȓ��N��jKg�;Y�e��2?E�㺐PFu!���BB�%Γ\����&5�K�wb?��=Q�A��Ѹ.$�Q]H���r!�`���#ھ���U�5Qz���D�Y�Z�gmjM��դ5Qz�ֵ:��b��o�]���m����M7ta06ܷ��.Ɗ�6�Ѕ�`�������ta0VܷK�.Ɗ����u1V�Zq�e�K�0.��y*�AO��"u��KJB�BB璅/�5$i�;~�rŇ��ya2���,��2�%��<����O�Ů�B�dS�-�~�s!��ri)x�N�#��a,���&�TOd�<J�y�P0\F�	e��P�]ާ���O�E�Ym��e���C�ϯ>,�b��Y��X,׋Ͷ۫��~ۙa���ɤ���%&�X�W�̴����ć1Q�&Ā؈	#iB�QLL5af�m�S�fCϩ�I�y�ɩM義�j&�M�@*�>�� 4�Orjj��4:ub���8��m*���ӛ<�2�1<�or���쬡�y5�)א��|a���Fl�2��^�^�9��n�0d�Fy�M��������=22��8wʈ�P���/L|G��!/X$<��w�'��Ľ�}g�#//38Y��"+�$�C�K#?�.��љy�F�*����|�d�$��R�&�6�lJK���oŻ�{iZ��
忕$e�?���O؟����eB�ə��;Ȯ�&9���,��G�����5sB�4� ��"�fN�t3'd�{3g`��d�d���&� �4/gd��3wo�Y: �d�o=��w���ibX��6!,L3� �V�|'�8�9<���q��"L@gi1C��d�h�F�֜�a��0����vd@��?8�J�Pλ�O�~��o8�m����9|sB��|s�}I�J�In���b�O����ݿ7eY�/����z�K�|����*�\��Յ`�nUti��­�6YC�Uѧ!c�*5da�V�;�0�p�ϥYC���V�,�!��s-C�n���!c��\��m!�'�}�'8Ps���͔��2�5�p�o�Ly �(8Rs���ϔ��2�35�p��My �)�Ss���єb>����)�Ss��xӔ��r�?5�p��GMy �)�Ss���Ք��r�?Ġ&�M!�c{�6s�ñ=5�n�b�	YCԱ�{���Hu Ff��#��1�p�Oda1�YCG�ԭ��Y���ȟ^<�2x���u@��,��{cz�V>  �k�1� o�p����@���!����%��c�d�^ x \�9�Hր����ۚc�d��x ��9�Hր��;��ۚc�d��x ��9�Hր�P5����1t+2Z�zH�z�i#��W0�a�e0��n��*��k��ڥ�P����c�j�U���Pcu[���������fy�_�_��O`�]����֦4��v�1T˯U�n|���gpx������hm.�Ã������EkD?,?��.Z���� �a�10?w����ˏ���_�a&���̰���%�x�e�������8̐��w9hѱ
�!C3T���#0C�f�ޡ�5DG%`��н�~�!:23l2o~������0C�f�ެ�5DG(`��P�Fk��R���z��Nc��0C�f��ƣ5D�)`��PU�5��O��PA�)�pt�f��UZCt�f��U�	ZCt�f��U�ZCt�f��U�ZCt�f�����PP@��-���1#):li.�e.i�a�t�T��~_mŴe������Z��ᚆX�ee��O�� �:��px�ȁ�>D?,?�J1ꗌ`��1�3I�~X~�`�x���:j��58ɱ�>DN,?��0ꇮ`��a�+Z�~X~�a�x���4Jè��#��/���a�i����A����(#Ѝ�Oc'�:�a�G��|�����t�B�Ú �����T�M �h�V�u*�& b4D,`�:�b 1��0C�J�	�ёJ�ac���厼�ZRt�f�S8F^��!:~3�)#/'��À����BAg��Q��N�y����P�p��ZC����t�B/˚ ������M �h�[�u
�& b4D�-`�:�c 1��0C�±	��q
��N��@���8�P�Rl FCt�2V�z�}.��'B�EY�I� ub�//+Ҡˢ�:V���Z1Q�k�C���
O�C�9�W��τ�$��9"��+B7�~R���'��~R������,���g���N����X)� �"�+������I�������{�Wrjob�z:{�#$��ނ��_����pY�	.��<)}�$�;~�|'+�l�{A�Ǣ(�K�� ���۳?7	�����y�p��l��I.�\Hk�7�/]߉�Tz�XD�W��G]��ljK��Юg�Z�6�^����a��@�?�H��*�&��m8���ͮ��j�f��j���[���Z��y��g{9|] Se&��|ix6��}ix�FZ��N�4<S�m/����LͶ�<���ƭE5{1�~�-<�ݗ;��d�m�f&F�;�5�S���6Ό�GL�/���t�6,�>����n��R8�!�I�
�d̔��H�<�r0�!�:f����4�?f�����ɼ0��I:x~J���g��G<w^����N�
5�M]�B�A8t~R���w��:�V�TF��p�=�	��YO�E��7A�4�:�[jz	�S��S&W��RפTWRyW�ϯ(��Ύ���#%\��H��:;R¨SGف��g�_�F���dE^*��n{�+�Y��j�F����*��>é�y��T�W=�UsՃ�\��W=���UO��*�wvq��sс�0.:P��[�����ƾ{e��PB6&��>=J�N�N۹�M����a�TN�M���#�F�ȱ1�<rF{���m��Mș̦��h�	Lؘ��+k�	ML��L���5��B�s�se�l�Q��f_�1_��$��f� ٩�a� o�cFc7yY�;��gzI|u�fs9*L�Z�(:n3�L��a#ߐ�QB�c`�!�0��]2�f�24���o��#C�}ӵi���;����(��&=^�FM༑	� �)�N�x�x@̶�v�l��b��(s}��O��*��J��n㿫�W/�~�.�q���!~8�ۇ��!�}�?�ۇ�á�}(<
ۇ�á�}(>�ۇ�á�u��`m9؝m=�Q��amE�Q֖�%amM�Q��EamU�Q֖�eam]�Q�օu�m]���p��KW����\���j��WY�D�d���I��A�9�#'N9gI�3��o���i�ډE��(�u�7*q��(y��I �˥�-�/�n��FXzEy���~p}q�/j,�+��Jo��
��y�i8u�w�EU_�!��ct�vv�ӽJg�R��j����RTy�w7k���S�n����Z�����::�z��nտ^�y�����������R^���������#y�����O��Nl�Y��J����}�܊���^2�f�.]ߖi��݊���f'J����٣�����ȹ�/7R�ocϿN�8���y���Q�~�B+��$�U�N{�G�p��)s��e�̒$�:�1߈�:�_-׻}��k Rv{~��.%JZ��Z�r�З�|%��ۘ��`$��ÿ�Qߑ�O�����|_��������Xn��]{מ���D������Gz?�cz�{2�����������Я`B>�5L���LÄ|v�o���r�ս��^�CS��Rm�%�� ��Zqߟ�qx�x�ǃ���ޑ���;YeN�J壘G��-x����G��&�`$�-c���\o�ʈ���*v5���%;4������,�'r�Lߍ��O�(8k�,�KL^7����욇,���̓?%A������Y�r�%~�\>��zN��0��ܓ�����m�T�˻�(sfMK��tՑ�z��DOv^�����݁P���{j����K~�9c��.��g��V�x�D�5��"�iB��0_FA�޹�~�OKY�r��V�{~�0/b^�i-ڸ��^�7-m���m��q�<��_�ɹ//�J_f�h�����f[�.�����2��r��]G��
��LyH'�]f�<����_� �q!�JHU4+a���XYI��znw�;;��;��?�=<�~���AsDAρ����Gzx=Pa�ףy?z���ب�Y�F���♒��/���t����څD������rZs97�{��> ��A��#��QYG�婺�^_���G��t5�0��f-���9�rDA���fU�����*������v?�}�����wWˢ��gYP�9�^�O_FmN�g���3���U{���j#�����V�꾬��|�pD�2��Z�Ä<���t�����cL�.�'IB�Ϗ��G�Ã�ͼ2O�,���l}s�?뜸��L� �<9�E��7��	�lJ/�<V_����k� ���|wt��+y�v�*Α�8�R��"\�lI��\愒o,���.�x�n�����>C��<�}C'��x��dy��<�Q���,;P�6;q�FDQ^&�t7*$�P�A��ȹ�d����O7���;�oi=}��O�;[W����oכ��y�G+9?�j��Q[���}����y�\��^��r�dE�e�Xd����ɊDj�Y�Ga^�v���yP�\�|\���f�:r�ꫀ3�S���]�Ӕ�n)o�4o�ڗc!d�ó�A���H�,���H<O�B>~�*���y�	iY6lay��������[�fo�.w3��z&~J�ݬĬ�wVn��ͭ����2OW��rb"�7r~����z��J�
��-X�b����T�Wg����f����r�v�+fw��/�z����˭H���k"��ﯳ�����>|�p��_˙ă�����Q���}�V�ĬX�nV���LNvfo�<��ۥ�+O/;���<݋���T��,݊�q
��TH��VN�D��;���{���f��;!*dǝT$����~YHE�I��r=����M�׸R�T�����H�>+,��9ty+��Y�qv#y��t�q��Y�ݼ����(¿���^�\�|�|'o�S9]*<O��R��&v׳��׏g�e.捻,��L�ޛ��潘��mg��*�[��˿H��Rr��ݪ)���`|�����?�g��_�\����oG�3�k�y�)�J���7�>_�[]<�~�����T7���:2[��=�'�g,��r�s��}��c��{|>��FNi�ͤ����r�f���W
w��h�y�AO[�Yl�H������u.��w��w��K�YY�]6�:z��ǫ�^����x�����7�1Z�g�|���ا?J�<�r�n�l�on�{չ�7o��;���UL$��z-����}'�������<�N�oo�ݯd��~r�k�/���g/����?�T����|����q>rܻ<>�=x o�����gQ9@i`ձS�7���l���~��?�TtS�m���/�������$t����C��}v�=�S�������s�y��2�n�/!������S�5�;�vu�W�{}գrf-G)�^�{�-v{հ��P�y卨�����l+m�rB�zԐTϒr�U��pUAt���7��{��e���t��Kq����/);�?�T������f�fB�C(��e�7�uw���;���L2;
,�Ƨ�dG�W�ؿr��
=R�~��FT��SI��O�V���s�hs��ٱ��yG���v�c�n�{i��˯��쒕��H<�J�����6��n�{�6��w����͇�w�-��Qu������7[:��w�̞���m7r?\x';�D�fS]�Wi�v�g�뛣R���{S9��fS�����mo�+�ë�� ��������~
����e)���c���z"Yș�G9�З���-�NΣ��Ҡφ�g���G�^��d��J��?��ۘPE�/5��F�W�g��Y"p��Bu�����uVG�]�|R����������9����߿<A�:�Wo��ƺɧ��U�D�7N�:�4���y�j��=(cf�eH�4hLMs�����[S�=�#�]��Hr����Ѿ�s���"��K{+6��P�_A��-eHQ=u���F������j�u1�Obp� ���=']ǣ�	t��a)���EZ����ޘgwv��^_w����]^�_f����o����#-�t����N��Őt����::��>-o��w�������N�5N�ѯ��-�1��Er<o A��Ɵ���<������t�㮚�5�Ïc��(�5�/��q��8�c�m�����
��2ϟ<V�=uP��o�7�}�����{���8s�su�'�?�*l����9��Cä���W��"U�*��.�����h�.��F�v闆�^8�;�;	�Y��ۛU�>��J���C���[�fMp�0��M��Ꮻ���jOq�!���B�ط"�{��ű��UNi�g��i�����Re��ݜ����>{�'_���ً7���xx�0:B�
oV����VU�?~���e��A��ˤ�(�؊Jכ�Ӽ���?����ɣgO�y�����=���/����v��=߳���ۓ�_<{>*���S�LoW�A��\o>P(�%��I���lw��r�{��?��������p[���{�m��a{�������k�lf��e}��[��'_�������hs����"U<;mC}��ϟ=�d�|n��fg6|gO�5M���i�ۿ�S���)e$�X͐.m���Mg���K�Б��DnZ��yƬ�!��i_�|���?_<<�E:��k�|��7��t���;Y>J���V�7���ٟ������-����4�rY�u.�pܕ��t@<5�1+���4Nz��U	ݪ�n�0u��T�ы�l#���N����z�Օ��!|ֶ�#]�ݽN��a���Q�;[�����"��bU�_������tz�>x}�_'��^�z�pR5��b��+$�jB�ͭ*༫	=ktV��V���A���i�V�:��Ϫ��:�r�kr��F,Ix�G��$L}��f��&!ɹ��D����(�U�y��Ue^��'���T��������t�C}+�Q�ڪ�}q�.��Η���t]��5۞�� �σyH:�e�l�w�q�uϣ B'KSUf$"'��QW�~��y���fIk���#��ӓ��Q�Κ��P�þ�����`Ф���]�wW<�;�?����L�r�W�6|2e�G�	w}������s�AO�!�\v��m.�ڍ~��ft��pEX�Y�D�ZM ����i\ƞeXҾ"�OIP��I�����Oc5�9k} �Ӓō��[�	���I<��Z�AM���n#��+�KjÐ�T_Uʟ���o���:>,��[� ��:<��VT��T�]'QTm��S���|�n��ŗw�M��S���o�⃪��/�Ny%MU��''_|�W3ny���W���z�ڡuQ���2]J��ަ^#�J�'���ld,�*ݿ��Q��Z��e�J�k)�l��o��V_?�9�E�{�`���aZ���[}�黫O��.����8�p|[�#=*�p|��sdkh8C��f�~�>��G̫�p�<m�]�ᰉG�*�p:�jNrq�o��ƭ������4��S�7��n��tY�V �E[Pٖ�i�,�v,o�˺���rрUQ�ĝΊ]X���)^�؊h����rPeC�1����(�M��i����..�����>�M�����*��g����3�P�Q��Q/!R��eE��\>ҭ6�V�׍��撺+���~d�8����_�0�k��V�Ӟ��)�z:�(f�h�i�����&�����}�`&L�'�d��m�vQ�^����G$?Nl���vOkt���z;�~ff��įlv��fx���-�dOl՚rwkY���Hc崹 m��qr�\@���1�ɞ�|�֪Z��U�0Yr�ze1w�'�ZR��^����.4t���
�t��4��E#qOfҟ�*�J�&;֌Bk���j�(&��k.N�~^� '����Q财�i��檅����7�L��-�n���0�[�VIOn�2�PF��N�㺷�&{�BnG��|�<�P3Kpf�C%P3C̡��)q#ʣ����WtSuj��U�/�,j�7UO�h8m7e�4��wM3�?gw�9�w:ϱsYMË�K��~�l�=�5��ժoPc�?<k��7�B�f�� �A��̠{h
��V݆�4�V��L��g`����{ڳ�щ�4�fuYo�gP�4�0�Ҫ;�0J�ѪǄ��I|GK��l4	̨����e�Չذ�b�k�o|9���NI4�;�1 b�hڶ���` �����h���X�8i�T{������f7�g�j��v�əc�mc�Y�X+��!�L#v��-4���q��Q.Mku43�Ċ �������M|+�Ah9lu�������i%z�ͺk��xB+�'�(0$�Z�8h�>�20�7T���,H�h�]>��7�3�F�5Ѽb���yr`�{��3��H]�������H$����r��M�'}�ߑU Ԅ�\����h�I���P�Y��Z�ن�H��l�cB���j���*�W��*���_�,����m��r���^�S�|��������|�X�������է�PK   ���X��g  n  /   images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.png�xUP�u��{�;�)�AZ����C�I)�-����8��P��+�{���tw��Μ93�pfv�,B��*�  ԠJ��&��q��un���j�	 0�����z�Hj/�w^z��^�V6 ___>GOk+7>W��S) ��AMI^�/�$���Ġu����������1�6�b���w ����(:��9�A�B`hz/�抉���T�K����%U�0�2!54����+|������#�lI�)���ŶE��V�c����m+�h�@.�����9UF�*o�@��Qt&��t�t�DA:2�L��K�H�e0�j8"0��h�����A�a��/�b�V�D�o��휞�H���l	}� }L�~���>��t����|f?�Y�����0)�){��`��o5����1�䩩��-��&�{�6�P��54v�J*c�?Ν/�yޣ���;_�����WF��� �z����ܻ���1)�?�n��9[��j��U�Ҫ|[;9�K:�D"�m�R����7 쟟[�ެ�68��<Sic�"�lM��ljn6b:m�&L��}�pj�������\����ֶJ�U5�tޢL���n�l�)�ox;nx�TY �J��y�I�@��y?E�ʯ���zZ�Ҍ�w�;��T)�?'Q�63�������W��:�@��e���4�R�I`��V��ʿ׋[��^��FS��'kc��������k����$C��7HY�T���H�"n���v+k)6���2�& �gg���;�>=�y������SAJP��f,����ׯZ�:஀[�?�q���Ǚ�UGtY
~s��^�F)O�\��Ý.�`{��3��b�$�[��H�:/7(���D��Y4�zV����;�r�w�Jtw��t��iYuI��>~ɺ��%�^4%����o}�͊��!b���k����PP�N�˺���y^�i���	?	�<��횇
���<疗9ϺN�s���Y�S�nF��r4J[���松>���]!faU����3�:ːG�q_�
���?�君���g��fٮ��v*�	���P�������)��Wic1�&��
�*�QB�#}�,���Jt��Ut6�c�Y�RY����m7�dgF����w�9f`z~���������4�)�n2~��m������遡`W���g'�x���!���+�y��Dx���/ǚ솎q��0�ط��S�<�+�/@� J��,jnn6�FB�YW�1�z���0i��,[����zUiQ;�D���ϽL���HN[��|o�����\m���UU����@�Q�������g�3Y@�/���Xޏ�w;�s�n�%߷�WtMfI�0�c�IUr�{��K�����a�u:S�a�n|�IY��ARĈՈ�:� ����;4�JMP�64���g �6\]a~��u��E��5M�e)����N;�Y���@̬�{V��ɫd}<,�� rp��!wL]ה��V��`�|��L&�E��LJSKy� ��V�;/�w#����(�.��o�L*��P�,���L��f���n*��/f����k�M��C�I��V�{��f�9��e��x�Wڜ{A���S�z�}������:L��3�DR���5s���l��x9�o!�b��9�!��9�����ӖJ#v�2w48SݷwӤ�Y��VL�kR��NX�I��w�L��/�����}��ͧ���^��hx��x��|Ԗ�+�鳵�	��H|:Cu��*Z��j?|8c�{�|N�1)���.LCCSu����L���(���(]�:��@-�/!�7�?�X��M�-�p�.Jjߺ$�s/ls͂��Eg��L�8�:�?���{t	)�|��V�~ܟ�����n��Lu	�gAOB�����Դ��>
�g���xԂ屙�WȖ ��#�!��{�8ğ]�7�F�G}^���8�xڎV+/��f�}�X��}�,�<cj{h,j���~f��gi��Z�陟�`�c@�3��8���`̂܇�7�7+R)wQ6����"z���:�*��F��7�|l���nI�o;u	%�_�ۛ�?>܃�Ѩ&~�	 ��:#K��6
n�F���4epftg��(���Қe��M�o�#�a��%�:$�O(���SH\'dn��DN�O�)�Y��"<����?c�Ǫ���	Y��;���ª;�lH(�)x[t"�"G��<��㬖�r®�k0�&�`��C.�"0��<e���a��@�^�c��",N<�s�9q x���f�\WOL�F����j�&l�f� �����0����=�����	�@L�6Y�Ed��Cy]���N��5?'?_���Y�q|N!u�ʜ�s��u�N`}���$~��g��^�z�qr	J^b�e�T���ouVT6 R �zynZ�e���ۅ(�0���ȗ�<Y�/�hm�K6`ϓ'�L4a4��{�щO����������"�M��8�;>������m+2/�O������2xS_:x���S���P��A$�޳�l�ϞY�(���5��l���M�'ק*������w�}�����Zq(㪯��ϣ�,�݄1��-����E�w�>�k�O��$ܗC�@x�j�]��O��'N�TY���"\���Q��K�iJ�y��1��欎|��q��b�ӽ�#W��T�Q��ݪ�6�E�#g}v�\|)&�Π��!��S�y���k��i�$��f�*����˫"T]P2 Ȧ��$-t8�j�QG �7��XV��#�{��L�v�&g|�|�;I�Q+>T�f�b�+��s.�	�]t�ۃ�cm]N�û8��z���׈0=XX���8l����=�]��x9��^$9�m��r��/���Ɗ(Nwn��X���Ea��z/�ejǫy&�G�A�1��u^�U���e�Rv��	A���L$��t���k󴊧b`�x�`�`m�c�[m|�q����%�`���tl&i��{CwC�W���v��3zB��/�0
�}���j�FχY�e��QeUNh/�e�违:����y��',�[`�Є���l�#�w�-ܳ�ע�yRx�DE�����.B��l<զ�	�b(Ι�O���5i�K��Վ���R�'C�2��Ut��v���R-�U���H��Sh��W�\h�a3Kf"!N�PyMlOB��	��ɦ��T~��p����&��.��`�|S�����YP�H9B��7���'67���!�2RT��l�K>P�����F۞)/���� y�I���I� ݺ�
혷7������v���4��YH��V~8�(�y�E�l#� ߄ϲ�̲�'7@�eV�M �:P�����D���U9&��*(h���p��`�V������Z��ڎ@����Wu���T�xhT� � �ɣ����w|��n�X����7��`���PI�l�� ���}�wd��.�Dj�z�P�1�sB���E�!w���Q�(�����z�Y���H��-S+����D�Gb1N;h	���4A���	��73o��Z/	[)*�PV�"6ӱ1S�$RϠV�+��_��A�>��2;DU�l��
r'F����m��;d�7V�+�YW�H����4��5K�/���z:©��/ؐ�O��n�w���f�eD��<}�?�Ҽ��_)��dz����"��Y(v�+cZ%,�`�UH��(4���ٯ�P�e�+�靑A*&�4Xf�%�#��#�(�C Tq�j�YSu*r.������K�<>5W179>G��gf^~�Xݹ��������.+Ը�.��� �	Y&Ic0mu�]��;LlV���ֆ]2a.�|�K�FE[o=�a4�X85�=�%�P����V/AK�Ndb$���
���(2�R��t�b������ޜ��R�~�kbs�ۦ�]�{��&S��Rk\B\c��#��o��x��cK�\ۖ�1̥܊ou��p�rZȠ�xu	焝��9ȟާ�F��|nG|Wo�bhp�Y��`��sb+����IK�h�=�6{Ǚ:_���������ߍ����B�"@sMGK:�`P�Q��Ls��A,p|��{'�ڤW�/D?EWp�c��؊�o9M��
��M�'�c�{y�z��e�#�F�l<�B��]O��%۰O%��<r�e5C�f_��!>�ν���g��_��/gL��f�#�EgN()-#\$�\�Y���DB>'d�f��d?���@4�7h�
ǉ9���x�5�������:V19q���WxQ $���%��56��	�2��ea$�E����Ғ	�tlRh��`	d-f�Ԓu���:&�h�S�3��я.˨��v�ٜ���j$cT��	�$7~U4��Βy���&��=���Y��!1b({�o��rz3Pǌ�:֦�<G4�R<E�e�̼螪oJ�e�=��{�ތG���#��Mx}I�����G���1[g���X��p��ѥ,ߋu�e�&N��<.Y�WNH�k�|c?��M�
�t>�,�s|�2#b��-j)�������o?�ǘ�}�U�ˉ�V.f^��q�`x�9��K�!m'�������7�-�QMs�E�`λ�_Nz3
?�;�e�͊��~�]T$r�Ɗ/U��
}B^���c�k���~���7�jF�.l�g��^pr�3��+q#��)������{�{�H��C���c�L鈈�B��\�c���ġ��q���jh���@d^�Ѯii{���;p��e}w9��l�����YT�'_!ߚ;���¥HfH�+�2k�5�ASF�j�ʙ·P:{���s��	��d	��pT��!i����x~p󂭡�RS�R\o�"V�XLq/	@�U`,0�������""����*܍u�P�xC�|A7K�e#,�b�m��:��*�8�NB�������X��[���J汁w?���h��09qװ��~�g�(�5�׭�F�J���_�J���b��5Ƹr����z:P^��kϹI��\��7��������%��|�SB�/�[Q��"��ƚrK��T��(�R��T#����-K3uwUi�4_I®g����x��t�S$/�������v�"'V��c���)ʮl�R�Fp�I�xrQ'f$��[������X�%Z)	��t7^�RƄ��g��:_�ޘ�K��������.���*�|�!���K��s�?��Rl9g����fr��F���f��J�CrVZ��_�S���!�Q�̛��D'~�A����W�E�pP!.QC~:�/�y��$�c��3��4��֋��ULM��W0Q�v#�C/�B�9��q�=�݄	 S���E���}�AX��a��*� WMa��ə�qOu���EDO��k�ء��NF"|V1r�>�R�ʨ+1�T��@	'��x-x��ˏ�g�ea�{&z��6=O5���p1c���X+���cQ9bǆ�����dj���[���d-*b|Hvցޫ��i�zeG	{i�*.�P�a*`��!���]}߷NM:V�hR��~�
�v$|�RP����(����'�c{!��8�[z��!p`�����B��۟�֚�-T7!��0 ���A�Ԑ��@�$�9	��#��AV��ZO�TL�����N���V��@�2�x�M`�w����@T�'��B|�T��)��J��o��))��9)ӢD��s�a�!8t��le�%?'B��p���?�F씿��������_6_=UbkN��Mj��Y�d�_|�{1D99k6��Z8AM��ƪ�����rF�Aq�� MWZ��m'FM����;-��<|��t�mN��a��O߰�O����O�',���;_�h��u���sm��$W�S�HĊ��ԅsv�wث
�� ��2E��4���a��y��ܖ���䒺���x���X�>/�X������w;Q��kG��J�ի�q �6ǰ=��I�u��F$���س]8���3�F�j��)�/!ݲr��Ք��4��l��hgf����c�&�IK��6�!�Q0���x=��]=���,��d� ������0;����=��i�@w����sk).�sOvA�y��W��oh��6#��Mbۍ	Fm�����F�F�2��PK   ���X�j�� 7q /   images/3afa6c98-60d7-4a37-9aec-be07fd386e0e.pngT|	8����R�$tN��J��%������&���-J�"KB�}(�JY��6c�!��G�I��g����*�5��y��~��}?zz[_���&&&6�׍��X?01�9||'�F_|:�����a�t����_�7-���>R��ku41�<�y�������=����%GW����������U&&!&��&���Kָ�ލ�)�N�>,ie�8z�ｰ�Q�>k���]��cr�c���e�kw1Cο�n�r�<��oL���G?[p��?t���7F��J ���}��)�u�������T���%�RtHQI�Ly��G"ovf�}��-��4(pTr�}�һYH�j$�A]�`��eE;�	��݅'�b%�ĦF�lt/�DP�����d�����sՍ�s���-�����/y �ȻX��e�g�П>�J��=H�m,T�k��kT]�t�K�H�`����k��R3�2�Y��O_�{��X��&�T���]U��+�^v�����sq0��96]�D�,潕�d ����6h�8��Z����-1�r���vsѱ��b0彄c�@��)��|�,Q����:��0�����o�t-O?�1�rͮĤ^h����#���M���@�g�p�F�(�J����pd��k=r��{ �zq��-MN[�]E�>Ò��!{��y,��3<��i8^j	G)�P���ʉ!!��[W�JՖ��N�����b���4|���N���.kK��t'w���$-���##��0ֽo��A�k��K�^/�u�w',T��}�E�	�i	��O� {���+m���.�����bmic��w��1��c+ۋay��؜=��H����:�޽[Y�^ȥ ����m�m�%{B��|F��=\��뚞vW[���.��h����?}n���ג+�KE��[l@ af� ��2_���X2�	�n����O�~����Ql���)v'A;1��7�}�Q&��&��#�d�^J�%�wxϩ�"Co���^3��ٮc�$�4b�K���#���e��ʴ�'z����f����7��f.o)��4�;�%]�'H��ĳXRˮ4�������3�q�H"��H�b�þ���BG����;���
��b(�}��De�0$��H��G��j �� ��C�*��X1��D�eE�@���]�,�m��*�$�QB�g�X�g@@���b�q����j�x�˂��ـM��BXep �r�t�ʉI���s�n6H��Xi�"I0��|,#�&��t4�/&wͲ��$�����Ǉ��T�iB�f)s����9�"��'����wB@#1�[�H�=�Ge���y���m��_7�:������ �����A�`a�O�eMS~����&��&^�N쀩ϻ�oʴ�D������$�(�Ѻ�CbC��<�t����G28�H䱹C�xK����� ��	���tw5��D�b<�ˏ����"_a�B� ��B��#�D����ŭ�~�~B�`�@|)�Y��r�L&gIϕw�57	��Z��(F��<W�g?�L���fz���؀g�]P�S��í"Fw�JLF%*R}ߤv�'��L@ri�%|\ǖ�pb�d$�i k�w1�T�Y*�,u*^��v����6C<	b0!ּ�"`K���7��C����Mlh$q��|�@�%6-"�k�OF�&�~�Mԙ]_�0Ҟ�Ԝձ�5���ќ���8vT��d��a%�8�r��3�N�Q\�Z�1:��N�䆸�B*�qx��P����t�@5?��_�0��*9�{R8�q�A����u��E�c�bJ��z�J��D�N�S.t����B�@�/�� �gh�[ [�H�����;R���So''�GqK[���51ӦT�/�����W�*4�k5���_a{H��^�(u��:!
-���Ƴ[
�,��Ä	�~X�aQu�~��p{<��S����*���詎?�A�-}ۯ4}	�S��bJq��pCLJLL�+)財E������[LA��VJ���D�Yb��������ހF{����A{d���������@������_��mQ�C�ԃ2$L��
�FZ��F���~M��q#�ā����׎�7�}�ۨ�ѕ�Q77�����mV�+�ҵqҡ����z��J�Oco�i\�ߐ��{�U�>�l��|��o��!t����������B8v "����>��jF��F]k�\�ʐf�c��1_����ٱ���K��I|���NG��1�JLn��/'�*�ˡ��5�-ڀ0r2={�,��)C����/$��v��^��������ׯ�n��x�����خ���kKۓ�N�Q͙�B��a�˟�CN>�z�Dlh\�C���nJ(Q��������6*:JNV�<g����5�Ԯ�x&�\� J�j�jltۿ��RS[�@"\k���+�Z�]i���GG��i�VG����s�V,a��F%�U˒0Bsl�!���U!;��Ш$����J����e��z�e'$�ܠP�U�Zo��jb��j�|��������9��N<#s������Yt�����B���҃Z�&�!,�(�<uj�c�8���b�ɦ���'���<:::87WXS#�@ԕ���/�?���N�����~jnǽX;f��}���	���Z�*	iދk�}��/w�r�T�����q�q%&JU/�M^��x��u�b\����QфYÄ����n���S鹈Y�Lmm-�P&+mث���x�-h�n/7%�!d(Og�q(v=��E��<AAL�ړ7�L/	v~`rw
~��ؽ
7ӵHaS-z���#�b�C�cw�%
�U�c���!����&�y EnH�GE�=�*�AA�^�sjR ��u\�0p��,E�b�v�-C���������������~�U��B���?ںfDd3��yz�*��k�QY��oPgnk�2o�	�)^k�f���:;�=�����?����	1�����];OI��5x\���������yډ��(�1ٶߔ:����,� �t�Q=|��ufu��a��]�L��/����jj9?~x�%�A��o�q�DL��=��Z�x_W�8'Q�2f	���`I��P����?��8����d#7�A�?nA �x�E���!el�%�4`/�����:�!���uZ���������ٶ�Д������D��z��g�4�l����q�Wf��?��bd�~�?؞�`��!;>В�l�1EX��`㤱��.pr>b�.�3ҵ�w�1���L^�e�h�t/�>����xezi8����KHioo��U�|09̤�T%>p�l�xk��S�#�ѣe�cɴ�6j�5+�����6k1��l!����D[�#+����=��O������C�Ш��}Lk��dMˆ�#�X���q��FN����9�Q��I���k-i�q$���1�s�q��%���2��\�6*�Z��.�%$@=�r޽����x��1_�@#�����..z�P! ��"�q,kD ��
���{��_�q_g�1�����S�@B����ܛ�Ǐ;�ʪ�Wt޸���!
ҧut(��9Kc8e7��3���Z)�f��;v��iK�{�4=�'zY����Kr��6��ntaI��c�y��?��Ib��acK�=z8��x/}^^^K+h��]S/S��7$��iIr�zE��5z����Ծ�h{���ݲZ�gDR��Ӹ1�?U33�3	����J����9���5���[��K$�Or����:�������Ȼ��H�U/�G�h'g�[ ��i�3�!,W�B�ϔ8�"�h4�=�y�c����o�)�F��fb r,��>��F�M�>�V�C�Ղ�"һ��؁��.�����8��9��h�hGק����9ɛ�2␋@�@��|\wղ�9ğH	1��l@e���Je��.~���{��)�2O;��x��n��9uXY����k��ɽ.���#��5�IW�+x!��,IP��߭׬�|�TC��~�-�а=�J/萭��7^�?^VF��F^Ώ�Y@9d@�S80�j[����̇�3H��mi*�Á�氄����/��k�t6�:¦+���k@q3����[R��:�����<=udd@�%I��ef�|DM�ۚ¹�R��TDSSȣ8���'��IR[��E�6�m����0M?����%�^�XX�#Lл<�ƔRP����O;8P��7��������m��t���w�l�^(��X�U�?)V.��@�U�c=ӊޛ��Г�I�e���m���:ꅎ�O����p�ף��*/�mi�tm�w���nsљ��OY�������x����F%��N�tw;� ��B��X8���>��K���j̵��M*Ss����+��%�.B*�3��	NM��E�C������|a������n�����m ߙ
��N���u�X�!ݒE��B���]����cZ1�=.1��jnW$�d�����[Ub��du/��(�"(Ky
�n�d8���ŏ?^���9���R-��fk:�q�Az1`3��6��L�Z��XrLa����r٫W����[� ��D��}}}n��Ds����k����R�4��vn��M>�<@}�6�4�"�~�'�z����/��OK��fwl[;G�X�H �"%5���@��K'q�*�z��K_��"�����3�+����N���*��Ռ�I����m���_��to���e;���M��
ViVV �.!110:��Hd��垆#��GC��X���X���^�/���O`2����Φ����*������D4�=��bDDc�-��ì��m����XjK�]i�}@\��=��O���S*�T-#Qu��(6��K����/ȩ_������Q�xߜ!KLbJ
bw���UW�
�����["��6[���x�!|�0gcs��@�/g���.)}��+^Xp��xbg3�9+�?��b[&&fy�r����9m�{刧�m�X�=���f�N������0����P=qw`�&�7S�GAyoO���9�FءBr#�	ai9*�PYY)86�>Y����N�q�]`���3�g)�c������x�n���R��PD��v��A���܁�>�UI	�� ̀,�Hl-{4|�(�c���lA�b���x�M�k�P������)H,,,�So���9�i�}����ـ
�C�g���a����E����vK�G���Ǿ�@�g�!��HW�R:�x7��� �R��sxb::������k�A�8�Z 
;,�ĂM		���_�/��5���i0�����UF6;�/���qAF����J�`H,TH7\�ۃ��d	�C���sU�T�Wj�R�(5�3d��g`p��c1�?Y�|}���E�@aF*j���NCخa;|r �DR���|.������"7�l]%����V3�l�]�M��\k�9��y�1��#���i)��j�%�\�Ç�pU�P��U0_׫�RW`U���#��{��M�FKWShC��f�H�x�_(Q#u�H�;��_~U�K���\" ���	eZ�\��c���0��ᶺ�3Z�����$:������8	T{�Jo��B��
��^����獋���Rrm�4M4S�h$A����
H�����/O4ѹ.:�����?�2�p��;'	+��@�~zU��5��~�r���#�.b'�A�j�>�>y�-����&^x�S*m�ɫ1�p(ۯ�2�l�3�q�o�Be�y�Q���2��ͩv���rpB�v�Y���[l'P��B�C>�{�St��.�-��!g�c�.	���!����73�OW�UlT���_��ڷ�G�ro���*�t�6V��p㳁�V�����-������_B^�MӬ��#�C#u"B�N-z�!�����w�[�0a�9t�r��l�RD��Pi����?|��g{\��WR$&7לJɣ�ベ~�D���\j��I�Ek�	�����FW����O�*⛮�nHnb��8���^��\J}��A�Cz�=q���	k�6��-x�#k[���MV~�F2��t�p��*>V�Ua4�ܮ���0-0���ߛ���ⳁf��0�p��6�mBl��q75c����M�V�o�X�v��hd@y^�U�;��)ymg��4g"m6��\���q4}u��\�V�Y:���l8q��򄲲rW$;��v1|���O"1���J(f;����ߙ�~6��E���ףX4K"��P���Ļ�d�ݫB��^؏��g�0���4a"1M�`{�`�qD5QO���:/����qqq')b]��u���H͉z�.��]�`o�-���ɲ�$�D��v��0�&O\�<K���FPc�G�C�bQY�e#u��Z�)�xq3�a�nue@<�>q$|�V�����]+-��W��a`���;*� ﶉ=��bY62b���geu���3̣�������+�ŋ�b/9WH��h��_���.�>�i�Z�brk�	{��qs%��3zz�;���˿�8} �d_�M4�����%
G� (���� L-��Ѷo���d��O5��b+�����I��֓�H��Q�B!��]�:1�ߟ����~o$�hs�͟uJ1�Yy&&Wr*Ի��Gr�f��D�Ի�:<����_�s�V��p^'�ב=rm3ǂ�cr	��{5o?�F�p�.r�R�@;YW�s[Wy#�T,}�x`��}*��%r�u����o�BWl}��+���%.y�;�ЫFE�;����N���>`7��z�B���K6���^t���y�Y��,i�s���w�r��A��I29dϖ�2'�50��P���< �$/��9F�xT&&�Y*��f�w(oa�' �oKL4z\���"�Y@C�����kmg��݉��:���bT��y�6X7�k���Vɋ�g�|~N{=�P�}f���Gc%q��@[[�+�C�U�k)�p�� �t���$��{7*1$�Q4��������x���+�|Pz\r�m*�>E>�w��X:�d�7i�3`�%�u�~�!k�^�Y7S7�RVL뒩��%�O~X2S �',Y��j1�*[`%��s�n]E}��5�pJ5��)��J��UBg�D�}q�gOA9��jp/���ID�r^<���F�H��l��'�r��+�&�RĿ�'dU�6&'��Y�\L>���NN��k�5�|�C#|��:�d�dP$1��L`~��<�Y��Q�e�NJ::�?y�U�ci>�<�N�u�tQ]c�l��§�3S��"����{��m�c>��ⓔwḑ��|��G�E�+Ĝ�l���(W��$�O��k��?�9:2��Ë�n��Q���!I���}~>'H:���URG[�\~�_�k�������!�	9.��XY= M	�!1y��x!T�L$7�����؛�>�%�k'&uc�����[%�K�~��ȑP�oT�H����1y����z�����'��eJ�4����Ѣ9��`w���7(�,��
��Y�)����k�Z����̍�-9�U����Hd���+�0 �#���`�0x�?k�4��.��I��u��e;}�d$=��u(��YZ@�_�{��kj�Y_9�� �?��o�D^�<J�V�s,v�l����I����Y�"p���u�G���_g�}��FA)�"p�Bi"�W��aX0P_>�����N}W0��kXrwT�)U��D �Ĵ�Ĥ��Gv����О�
��B:<<���kIz,��r����c錪��+��͆ʞ~��o�i4`S��~c�S�.�fj��^:�P<���<��pn[_k��|�U�K��:�(tؤ���b��	���D��p���{Z�p_��+��Q���Q���u�M�D�#��PW �Ĩ�w \V�D���� �c~\B�RA�R�J�YA
��E
�i�^y?d�⶯���A�oҏ�/�C ��.4c��JM�J_��-2�5&�S��T���퇿�ª84�=D_��ec+!�P#���;Os畁FMP�{�ʼ���hVE&���������+���FF��+�M�[�9��`�k6���cY���[�	�>n�c��G��}�ޘ�H![kW0���Oց/rNV�� )�����̐�֠}�*L_���?-���E�~������y�u5�Ǣ��$N��T���m©I�{K[�B��-0���/���{6����@��%�c�6bB�c���Q_�Y�{,���$��+u�gu<@�gǑ�Y�����c �V\c.��Z�7n���}G[�D�}Y	[�������|5�����Z[Ƌ�\E@}�IY�?@�}s��&F�#�r2�H�U��=!����z��򍓗<Eô�N�\�����.��"���Ȕ{�s��L(7�S���ؠ��?�Ϊ70=�u��#T��ЄWTp^���;��b����c�Y��-��	��̠���h�١-{$��KtS�Te���1��$
��:�"�%==l � �F)����J
}�b��_�]��z$�޷LG[��)�� ���{�Ѿ �����o�=N�b�. uۃ��O�k�Cpp'DiQV}���,����Μ	���PH^�G�e5���4N%&N�eY`�M�� ���8*�� ��'{�c�"��7p��$|ڸ&��2�C�C�l�G%��x\~'a& �ݓ c��ߛ�w�B>���x���bv�9��u�����;�^c$x�om�ɍ(?�5�5�@sUUUy�M��gD
���VZB�)���B4 .}���5�4g<�np@���α�@�7^�m������}��κʘD��2���+�u%�E2���A��bA�M���x&��2m�����A16�[P�����+;�]�Hu��u�}BK�t�9Zm5�$���<Q����@W ��_H�)N`���R�Q���	���A�!��f�/<�Ϥ��GEEɪ\�}�z���d�r�W��x]�ɬP^^8%��@��� ��_�| |�t��)�x�z,�^����,���~=�o8��H$Y�ښ�!H��ޕ���,3�~�(��#.>�r}���O�^�5ꗉ���Rfy����.V���p��k.@����γz�֝>Q��ת��jq�F�C�]1�IɅ�.�#�O��+��C�)ej��gR9���ҒS�/-u�;i>-W��[���~��m��
[��BR�ɨ)]�c���j?��N��/���<��Cl��L �����$~W�t�hеV0yc���,�`��i�� �y\4(����q^A<���᮪[WܰߞI�m��Mx�����S�z�Ma���n����<�h>Ax�٩m]�^΅�x!}��)������tB�>[��o���w�)�o+�l8�@^b����Y#��p8�8tŗ;J=S��C����e����Y9�R�>\���י^$'�S�n뀹Sz�nq%s���XW�S��x���(��|?Sc�V�i
����'�'��4����$|����giNO�-�e����f?b����� �=�q�V�����K�q �D�����!�§/��������g���:;|�^�r�p���d�#�2)|\ܪ?�k�p�0}�x�]���i+Pպa;�j�/�n��ST�q�u�iC����ދW��m<�S�8 ��b��ղ����=�I3���u��kYx'zk�#3.�u�E/S����Ew��xxy1�?�w��y9i��d���[e9�lV4����ւ�SMC���U�,�c	�`,!t�d�ᮧػa	�7�r�zU�vv��פ�������t�@��d	�Q��ge
37�d.&��:��GP�����_���������Y���E
���m�k�;�x�r'MS�kn�Qu��A��^�Ҡ��������_�׎��C�[�z43t׺�BeC�9�����yTܗf�ʱD���iy�qBxo-��{��M����+���(�W�M���FkW����Me�>��e.��1C� 3�#Z-�G�Xt2i�F�%C(!W�EX��#j������OK�ǒ?0�7t������H�Chm9bO7�^��
l���9��n&~�����Ŷ�_w=[T9_Rt��D��	�R^^�rQ2�X��c�E"S�d��_����w�r��r��9B�A��D����6�Ča@���"KE�=���F��0]F�,p�y��f���Eݛ����_1��c֏�" -�)ht���9���\X��e��w���Ӝ>������B�*S9p���
��.GL�<�@��=�ֱ�/ҏ2�DbB��n���V�Fd�������?��F�D-|�`q��x��c
���[ȃ2f�i��]ڗ6JNK�]�[|��viuB9pj��)88�21L|L���<U!C}U��Ω���~DI�
9�JZ敻�nk"?i�u�.�k��z�����^ʞ��l*�`�qm/��LK �����7�߄�?{�������������O;��b<����.?@ �^��P' k�ڹ�zF�4j��A4oЏ�t��RZW���!Сx���I�XЬ��,������K����ʆ�7zՋ�V;`{�A� �ݜl?R���H�_f����ـ�2�X�зH֓[��n��6��ϸn ��u��S0�c�WU0��)�n�'E,��]��]W�h��6�;�zh��dT�������,�C��e���lޑS7TBˈ�O�H�g(��j�r�d�?>����r���'���>&�Xi���ݱ@1���o��,*3�ѕl*���G��������p�{�Bd����5��9$	�|!s�u�VU�03�n��|�}�D�ggI�6�_��e���A=>	2���ze�g����ۤ͝����/rS�M��$���V]Y��;ԡviu�:M{^�k�Lc��a��d���1�ßΜ�A'���ڢ�{����$�hB�:�/u���@���� ��O�"}���ݤޒ��|�X��I�ORA敘k�t�^���V�Jo�t�$��Ҭl�L�bA�Jd?���5E�QH���:�����:�Ҝx ��s��øW��ᣔy!���{�U�h��\Z
�O�����OR�����h�,(p���v>S�O�����8z�pU�����hW����B��C9�"�I�w��3\W3��v[�Q���NM��yv���#:LC}�w��v�m��o8�bMB|��+\�e�̲�IS�?
�mZ�� vOf�&��Hj��-=G]���RQݣD�*v�]m�h;�]�IT�;�9�Jt}Lo~����Ӷ|n�z�Hjn��'�<���?�Z���*�wֱ�`����������s��i{�o���Q���9��>�Y$fe�v��������7�_��� *]kL���I_�mh~��k$nk�o��-���@r���o����z�����nb F*�l�S�̘�z����""��	5��5Y��㣣�A������b�]{��9Z|5��=-}&����a������@]����=��M�lt�����{o"������	�+�X�#1Wj�^��KH�P��}���>?!�7�	���f�Ny%Q>F��\@P5{�0?�����ڥ�@�4�d��Y���52�����Zn�;t�7��q�ӯt����x�+��x��kBR�bO�r��p�m��&�j���V���&6��3�,�~��p�OE���@'6�d������˶����έ3zz0�yi99��j�a�\���V�r'2@BR�\&��s?SSS'W׾�9����1����a��
h���)t҅��x{��i�P�؀faW>�^E���[��3��0���;�)�8�o�~7�O��о �|
�����x�l���,g�����P�|�i� �i�u�wR�X�A���!�D������Uν!�G[94_np�@ y�|���0�\5�����Xh���D�܃�uW
]U�߾e�͑�Fp��N���k>O(�y�~-(��ƹ��q���c��i:��#����&�sE~�Ĉz"oP�S��q�Z`m�ͱ�����������"� X.,��Դ`.����j8��Z%.���^�����m�,��\R��X�؝�B������NV���͝O�$U޳�����4��W�83��_ۊ܎�<����ӽ1�#'ǑJ2>Z��<�-����|j��<jG��ER1~C���ڔ�m�Z��>ɂ�[�pQv�1�e�D���Y'W�N��&�_�rq��]Q��u���O?�?�a��/�rlt��
�0��k��z�+Es��
���!JI�A�	���c��qrjj3���n<�@/�==8H_)��&�p�&�V�&��r�������F�
��k�v
�pB��T� �� ӊ��VYxdhp0Yr#������4�����]a�����
LqIIߋ���ѯ��uzKAΜV�j��
�I�����w��9M�
S�$S�,��_1�t.S'������T�֐�^�z������	����������+�[ih��Պ0��j6��2����D��!PM�����g��YS���EXZ�������'�5����gh�,�{�|Ҁ�xW�^��4孤����D_٬�Ԣ{�n
��^zNkZ�ƫf�/RBqY��/�/c�h��z��v�tW�������Q���WRZZ��V�0�ox�����E�֪�a��^�����\Ta�V�G>��Ê��YDݶ�7�U�f����..�箮
���7��j�s��k�z����, w5KNV��4a�l���蓶�'4�1oŻ>T����� ����Q_..Z��?R��{�SsϋSs����TيV�����'�@`��rd��D�\�����S�V�+���2s9U��x��(�����F鹽n/�A��!:FfZ6��s��q�g/*�a��������;(������H�ڔ��F*)5�х&�E{���ZYZ�#�g�_e}���Њ��R�����&{��\F%��z��J9��ck\||}:^@D%F��p��[Ѐ���Hs�����Q��n�ȣ��ô�5���q>���[)�R�#u+/e�q��Dt�>v�Xz���F�}	n���hɴi#,��Ʋy9��C���?�ySW�7�57���1����3�� �<	Xk6���hA0ƇE��DZ��3�0#O� ~Q�8=�_�bt�>�v�ADMM��+Ǟ�[K?�۵���UD� ��9H�k�W}����(���Y�ؠ�����	Y��~z�Y��\�*��"���jԡL#@�;��G�'uΣ�3�S���U������L,,^���a�J��� �����<~|��TS���VF�ݘo�G�ƚ�z���jߣ�	��M`��Z���DJ;��S���+(�U���ߚ9��My#u 1�G���))��UTT���t�X���}��_E��x> �<f�͇of��[���ײ�Fge[| vD$F�'������R��hv�De �u�x�j���j�j�:�boP�.ij��ϴv�B�E�)S�����{L��b?��x�GM+Ԃн�V"�੹{+A�����"�9�Xi�W~�������Z���9e��2@"@�9=��B��$2�}�qYÔǣ�.���yV:�ޟx(�d�.
�nM���(ef�Bh����.,�|�g�ں&��#cK���bqu�V�N��\��gqql 2�@'��[J�u�HN..��<<�I�}��Y���U\�F{�K��[��w�T�܃�s��l]I2O�W$D ������τ�Xmd���ˏX�v�M6t)%WD��]�:���� �ޗ��D�J�5�#w��ź�{�j�S���.�ړ���*�&�u,,F����"y��M|�N�`P���8�a��jPq����-(r�Z���Ļ��TaC##��{�]X�|}�0��;ø��� �<���[*�����<�0%��P���:�S��^�;_��������ȲT�Do����V�ogUz�A[RRn��!�hx4�Q�N�β�Zh]��| �X8��C�moz�{���h����k����������#�éiy'33󟫤�H�4U0��޶���P�|�}Krs�,�M��-��T|�b�U�	��B��.֞��Q�!�l���1���T���eJ�v�>��KL��W?�KH8:9�k��dikk@E��%`<�^�-o��@7T���m����έ~N�C�zQ�X��}�N�Z^����8&&�`��u���p%u��ř�}Ch��2[����o�JJ�'�^���7�#����>y�(��U]���X����1���j+xOD�+@��G!C:�����񹦔���"�NN>�W&$q�W�W'�:;���"��9;��Ղ�=��گ8<�Ijp����N��qJ���H��&$o*4�0Etq1���&A��W�ׂ�N���2�N��漇��_W��U�9Sz�ӧ�~.���ލAl_NE��s!3��R�>��|LaQ!g���HХ}�P7�A���`���1KP�\ �����,�j|־�m_�";����C&�0�����}����T´,"������^7.xF#A@m�@����G2%��
��˯�٨�h���=+�W��x �����%���(y�`UxI�E�[�����h�k�R5XYYY\P̮W��������� l��,�~5�{�_��Ƞ��_�ȠJW����x���]��ߙ�lӥ�k5�,!��Ԥw�j��1-fqU-{;����7�o��,R��ŋ��mT�,�f�Wh�M'V5S������\���MRG��95MGP��*�J�-\��ÁޖII��3�{w�Q�oջ�B)��"-99�6��%PC�b�r�2I�@
��|�@s&�G�/���1O�}!uT��(;��jPD`~��[M��g8�u)��?E�X���yg����y�Pٽ�v����A�T�:b}&���A{mmm�Y�i:�����pXk[G����H���`��� g.���[7�yy������gZ///�e=1�T����|���=�K:���mР�Q0����{�5��.+M��-&�@Rw�݉�)�ʄ���w3�d�DvRO5p���th���Uh�d��xys4��M��\>�f��?<\�]��Y�k�P���i��!�����|�}H��S�x�%��_�~y�M0���Ϯx�zp�8�M�7o�� ��L@?�x`�ϠEx N4�I`|��bȫ :%*E�M=�a��Ӷ
'-�dz����@�H?�����Ĭ�]4@�����V�A{��b|Б�jAw���;io0��x��ҷʩ}��ā��I���=-������;+ |ՙp,B����'Yގ� ���hwu�Q+´P�=�����{rRc�C�j�j+M�X�����T�k]`}>DJ�r
Qo�� 4�?O�'�խ9㶴����n�o@��^s�j{�rek�3�*���eJL�@�=ff153K�f�__��d[��1g���ރ��hW<�,��e��0(��^��_�RR��2��bb���������i��^l�XR�0�ｮv�rY�W
���	����xjb�E�����DJs���vM��S�KG`��h�/�5\Qv�j��UQ�s�W/�&s����$��׵h��ۖ1��j-#ݮ�Cn;n���xA�,?>|�I�~Q��q�$B.Rq�|��~���k({�^i|���)dė����h� ��C}�u�dŚ1��fbfZ�=3��~EC`�����P�3��D{H7Qǲ��u�Г�.��Bh��zj��h�o02�4O�3��pGgg��Ӑ�.Ӡ>�sc
`�.����h��ϾރBͯ<�)���A�*��9�'k�<�rm�:�DҀ�q�ݑ�t�pv(+-��r�$m˝<��m�=�{cN�(�f�/��@��wH`�W)�KI���+p}E�Q���r�j�R=�ԤfL]fpF��ݏ��0�_���ms �4���������1V�z��k~�qm��`�Y[g��R���r�t�E5`���K�9,D��*���n5֌ޤ�`ٝ�u�Α Y�=85�3]\]�%�e�����V谬�tE_�kKkk=�\UF��%@b�44hQ�["��Q�����ktx�#]��D��J%������ft���)'u5��+�|�WRRb��w��k���`W���I�fcph~-�����������MM���"�����&���
9���Pq�E-� vܻ@�}�zj������l�+� 3͝+��;)ꚺ���U ��*��C�
�|�d����B����~CqH�mi0�U^__:S?�+P�c#����s@� X(F��>�_O���$�}T������}/������@ې���lK+��#�5�e���)���^`	+�P��>�ޛ��
�S��\̲��Lo���T��iq��)�� ����X��6���"7�a��,��b�R��?�Z�:|ʹ�e��;)Ė;�ַ͑bc#h�|&�|}}��|��¯�b�\b�/Ў9��EL��צl(�ͣꗁҚ�a��B�7�aU���@ �$�/t�4��K:��m�pv�1���0f.5+�]����w��?�{�PTLl�qD��d��� ~.��:��,m��&?]�P�+t*���ҫ���-qҥ������r(�fߪ�x���_�~��9�Ƒ�h��>>���0>�����i���]Ɯ��ۡ{�������LR
����t��JGlV��#v��*������X@;(c�;вK�2��MǬ�5�Tr�07d����.zP����"eTY	���r$��(ϥ���={�U���>0
��C�/6�QaO?8�[�#�I7j��{U,-ο�V�_{.�lLfu�L�q��ʺ�]D�a�[q]������z�t�������au���e�t��+��jVaTM�"�N;��* �5�@���m���� ����I�WB1Z����|cj�)f�i7DN^�\f������+������冄\5�n�n=���I� ܞ���CQ��R��|�	�$G�s��0q�4��L#��qqq�++�^����ј�*���VS���F������gttל��D`�۽H\����N���H�==�C�%$$�Ӳ�l���N�.E"��|�{���.Ćª�o�;Xc���7&�6li���Ӕz@髀#�vpo(r�>�174�p�2��)j83�tt�4�T&<bH�\UY��`�x��@s�_�ퟙ����q�l� *��ފ�����MQa��Q���8�q5K �P�,��\�s�1����;>�q�/��m\��4�W ihh�'W��w���Ѷdic���������]���oK}��˺
�p�%���H�����+ `�ެr����**� ��/�QӃ��*#�1��5+ P��^c��Xh�Z��V(��߾� 겖^�g�_GT,���|}z�fhS��"�ଘƱGޛ�����t�ɋ�PYi��i]墼��|�b�x�2�<=+Km�4r��D$S��8űwZ]��-�����(�!^C��Յ��r�c�[x�j�C17�]�1䴗��m�/ի� b*���O�u�lG�5v'�9�y�����d�rs�?��t�>�Ӳ��oSX5?b���4���Ǐ�6�~���tn/�5k�;1RNkc"v��fKϝ��ȶ٪7K�,=}d�����W��`����^tIq�m[��>>^���b�X7��m5�R�!�yx�������f!;Z;��SWA*���w��/���ŃSX���͎�>~77��70	��x����B�\��7Z�&B����=��J��aT� TTwU�"��D:�T�U�"�UJ@QpE�ҥ)R#-HJ�H�  RB� B������=�9����3�<ϧ�̝��9���V����i
z� rO�X�~f~���p����w�;���acN�I�������l���ٻ��<��H��cd�����o�ÌM}�����]M��h�۷����X,/\�|c�������>�uwF�7nN/-���I��>@K�ֺ�G��`^�20X�? ���<q����o��"��{/��P֍�:�D�,>����j[X�>}�I0	{`e��|����ۡ�*$IX�ms����ݾ�h�����(erwsb��q���%�m���ħ[�:���6��Hľ�H�������$ܗ���&�]QV��ؑ��V�P*p��w��k�r0�ި�?�w��Ӹ7ο��k�-��4�R�5��:��؃��	Q�����V�N�T��U{ͬ��/���#0^c^f�O��~Ak��uy���a����7e�ȯ����XH7a.J�pG�#g\ϐ��(�����6�����O9:;�J�Wp�5iNO�(ݛ,P"�<Q�����[�%<:.��Y~~����m111	��b^~���y�zx���t�&������X��<Y�7��mT]z�a.*Woz�!����:��`�G)��2O����w9�o��t�J9[�]$v������T�ؕ
����(���`T�|��� ��,z�dR��Vu[\�����n�~���Bi�Ww۴��cR�����DcӀ d��%�O-T"���iP#=h��X�G(Ƚ�p*�4ePZDMi
�ˌi�a$��|���9������X"�%�H��I}3��(�]4>nc�u�gfF�>}  (��O�@)�W���OTA[�eWKJ���
�l��1H��_�!lRâfm�ߤ�پPߑ�6WW�Qw=ټ{~^_]C�� [3�y��֖d��o�"��ȧ��	9<|(E5#��Ln،c�$ew�K�:�,{&t�"��Ǜ6S%��4Zk�fY&�W��x�ӡR��!s��Z��hm$5�$n��A�l]���r��3)p
��|���c��7��u��G,�P5�y�8�Y.�����
�<�b��
@{��| ���+G��}���h� E�
W!k1;`�|�w ;���b���O����_�Ii�Fӗf ����h�������Z��%���[�.��嵬����gT���q^cMː��.$��.�k�v�NN�˂��y��<�j!���y�SJ﫨�
Wr�HL���/�n��M���C�E-yy��Z�4��9�/��'!I�J���r7���\!��V��ޮڊ�YX`K;��@��AN�S�r_/����?�1i�!�9ﷷ/�~T�C??U�F�W}T��VE��Ң�`��Hr���JuH^�{�7�[ec4=K%ư!y���!8{{{��R�;��O�[�c��@.)Oe���{^��fL�I�a��U�&#Eރv3@�h�!0��ɹ��|j���gf"m~[�(�u��S	�9'�h��\d�7T��-�}MH�P]٥�� HBS��d���߂��Fv��?:
�.��rf�K}_.����ގ��xy{;�;Rf�q]�,.�/LT�v@���&�2oqѩ_�{�DE�-|�4楮�jR��h���P�{[w�����I#���Q�*��J��ȍo�7�DiS|���EA�~ve565U�!�1�]V��f����~��2{�Fä,��{<����>B�g��W���v� ��mַE�- ���E�JYȺ �e7����T�.�Tٿ�76.n��#и�mN�!�W럤l��g�y�\Kk��H��|K��wS��2��<�>%.��U����t��p~���J ��յ����70Kg.��ދ4��"0"4��T*�[ӂ��5���0�P��+�R0~s�g˪���8�8��fU�V�p@�.|jM=Y��)N#E*kb"6S�C(ܳ2;w����s��@Y�Cc{����0���HaLt�k�����ꩧ�,HaA� X��_ė���\�IX#��"31��_J��Y�5L.xK�,n7�(��a�\ʮ����0K�������"Wr�Z�����{fU��l��w����D �r��Sp9�����m��V��!^��9�l����OI���4�5��˦���P�����&���d�����_�Z����<G7/TyR����Y�U�ۜ���We��4��(�a������Ll���"�fUQ�E����Ռ#�f�c���w� 1jd��~?(��I�HR��݈��Z��]|P;�kə�.@�I�:��WĀ8ڻ�/��37�N�2#�ڿ����b��$�nD.w,��6�J��;���#s������gf^����{a�
��G]�>�F��X��������}-G2�ʓ叛
~e�� ��#������e!ڴ��I�IL�QBOV뙘�|e/���	�/�jjX�;�qyV���ׯ��)���׼�~���wrh����B3��I�^BCG���19���LP�7'Bڎ��Z0T7W����>C�Z�쵢�N�L�7YG��:��\*9�^ZT�Owe_�4�3`�u������J�d2�Ex�J�T;dw��i.|`�@�����޿ln���d�.uW���t�?R�,,6Nݖ�!�$0��	��d��4f�
���{��-t�*P3V��>��/T��ۛ8�\�pe-��w�F]]�K��K�.9>|hz��u %#�U*���цz�K�
�z��c�ӄ������u,�N1�2����>H3�oG��8��e
MM0h�]�2��������(>�� CL���Ư9n�ŢS�UO��N^ɪ����^����s@��}H�ԗ��KE��{�B�Z詳bs�2���%ҋ�b��3�����\���}��B<��_׍��Ō�g~j��@���&w�hС���(�8�w��w��5L����6ȳtIj�� >>>�����P���paaa^z�v�'�� �)G[?��u"�<��T�H�e`��8�Pݮ?�H��6g��NǢ4c�����2�*Ȟ�۫o���"R�.J�~�%xwh�hHp=H�4N���ʳ����+��W�0v����{��*pL��ϗC�U�2=m�7�嬾��!�K<D�2�韮�
�{�x�H"P�ԥx����(����5�ӡ�ɀ(�@��XX���b��?#6/EC�'����L�&���E02m�����QZ��A&�s��Z�72Ҷ��2%�Kv�tt���SL{=�d%�o��Y��1�{�Ҕ�r�1W�b�k`Z��j� @%-}�H|�ߥx|�u ����������]����������L�A��W��RY�������/�G����,,�.�4�l�6��:��;�7�2���^�]
Hg�?`��m��I��z���bm!n[Ǉ6�"1v��_���#o_�Jn���/��I���՘)�BⰞ+ҩ�>y]���[�
��7>ߘ�n�e7�;b �ꔟ���a��h��I�I���F0ɳI�3�Tt��퟽ v�ֱ@�s����%�����>��v�j��N\�A�$�� G��](?e}��wg�%jcw�3�	'u{���N���@���+��6Y��^��X��ep/��X�Ԫ�E�x�O��V�M��SP14�50ԩ�<">����<{���dE]���}9����-�����`�8ϦDP�I7'���g�0��t#7~́�r��_���P�M	�V 	�ChRQ�7����?�*�I��S�d��쒰
o�U�oF� ջ<Q����uK��(�'�	��4��2Z�ڗV�)�v�Qԅ�������iC���[�f����e`e�-�c���;m�{�[���*	���������)U8DZʰ*�sH�D_9�g�跽~�k~�/�o{���4�/����y��-AYB;qnſ:!њ��q�&�]�c.�h�$�̼�rX�&#mCp�=x��?V5Gmz{/��}~~�Q��������8��X�� 5hc5�������
>7K"&y�6�����n�U��n����Rxe�1�����Ǒc��"���������|�q�x������b��(+ ͫ�a��566u�8���w%Y���7W���q��3�$��>��X{	pߕ����or���,��éd�.�����=0y���&���76�f��-&W'__#]ݨ���R=5TR��d�l���I�����jX1r~�(3%���b��9�,� ���"��Y����n�Z�_�}�N��f��tH��MOgꪶLʮ���*g�a�e�=���}�$P��B@	w�����#�� 	M���<+��/b��CջE�$%F@����CV|{p���ԭ?W� �kt��Z!�`��;x/˿&�R�x�k9������7<g~6:S�O�5h>�vFD�������y/cY�N��0γw[D���_q�:�kCZ���TwS�*�R�d��o[�ޱ(c�j=
��j�2�^<*�hJ�u����1��mm��5�p��H@��6�4[�����a����5���"��G!�Ɲ���6��2�*�
��?��*������o}���iM��%?�x��6�^�V����)�H+�{q�.�v�:�C�����~	�����^���x�UV5+���}:\�:T�9IF�����l�d��|~D��:4�r�ad;�腽`�q��~�(����P])��Ex�=�V��(v�5�~��	�,��f�*_�l�u�L�P�O��@O�� �D�E�t��	�$h?��x�Ω쾤QE�	�������R a\'S&)!g���R.ƒ��ln� b[��i��'��C.���i1�������&��k�W7NPF�
���z�
�TV�Ju9e�w�T��L�#g���ي� �Og��ȭ+�`�'ɏ̀����1�<S�|(~}C�d�~�~bN(��oM_?|�]h���dޱ����tV��x��(�=�_��0(���Ac�j�dJ�7d��]hi�!D��Oٝ'��u~����/g��ů0:�v�*�����"��
E6��;B���v���?*��QwX��)���b+^k����5�w�>�&ppk��_�J�d�*9W�%kP�w�9�?)�A�����b4r&�`�r�����h�!�t.�~[ZUQ
z�N9nv�g�����Y�$"��w�,S����s�$���@��w,��׫��)�2,I+~���(K�*��'���5%N�r	����AN,���.��_9#�j�;�v�bh�xJq�ᆠ����L �z =�c��E�T"H�k@(Xrl��}���O��Y��Ā�4{ '".
t.Mu�#�ʋnkk�1A�ÍJ�s���YC"Q(�ԝA�ӡ<���X���d2f���	Q9�#P�����D��qȳ%GM�����Kx�Q����7WO5�C���$J��mx8+�����w��!y�o�T�n0��6<-r�Z���~y7�� T8$+K�6�+����93�N��T��Z+�:b��F��mϛί�x��5����|����ו��?ip�wg?wx��c+y��ƽ�W��z�t�]��O���
3��Yf����_n��*�b[)�����"�E�U�;�"�D��5�������ɴ}3�0�7�s�����k��]�	�X��Ώq;��7(|J�6F�"��y��dd;��#k�'p�n��M��w��+Y���)ځ���;�4j����#�].���/݄�$U	U��3�,z�vic8�E��_��*��A��&e�Y7) C�x����}�z���sٞ�����bblj�~��"�[��g���o�-��YYY�R�(��`�	��/_�(݉���5
o�cƜ
�v1V{8e����3�y��������ó�����
��%����O��-/��-��$bN��t�� 
�t��s��D]B�Ѝs2h	����U�>yBN��� ��Bq��)�t����"��qBC�hu�iu�Nn�'|�S��F��=>������l���
Z��HJJ�(Q���~��+��[�q���3���V`8ۄY�\�S���&���A��}�h%Z��l���'�>}�7�$�2�n��1�h+2��%N�4*]=?�������:���w�(U#gy0����sH/Ѳ�omC����	�.m�3n�պ{*.(��n"���=��Z�~@�1�peQ㳍��F�U��t��9�,9��SA
t�8ŗ��##i�I���aFg�F��L{�������Uj1�"��ǳK�=4]fs~�֯!v��P�F��6��;W(���v�Ͻ�jЄ�0��s���,%p¨7���>ʱ<ϰȬwaA�O_:��|��F������5�vJ��5e����]5�Ϗ���5���J������v�����m�N	�0����G��GiiU��iߔ�?�/S���Z����ro{�r���me(:����;�Z9���Ռ����蝜��;;�pG�GF�$f�҂v��<h���!������E��[������(«a/ �CB%��f� ����ac���Τ@�C���(Ƨ����� M�W-���_��^P�L��X�����Ӯ4�حO��9BEo���d���������?�X����A�BCò�ڡ�Kk�����}��l0�QD;E������x�L����־}���3/3�i5����m������!�
��+��SN��5.�gy�y��q���X���-�(����G:M�[�h�/�3h�#[�:
t"��Z5?��x2�Y���ꤢ�{���Kp�yu,nWd�B�8-��C�٪x�;�M��#	�.b���5r�%z����;�lyiiԟ$`jyǷ!F�9i��&yr@�t��g�R�N���Omй�b/�Ϡ�R��"�.,z-N���U�O8	�V �a�©^�
�>�ڍ��>(�V��%;�75@5g������!0�U~�61���8��u?�lw��.ޔ��`��h��di�
�63��1X/.6��{�� u���w/}�7�<���k�����S����*iG#���A��T�=y��јV�ڍ�>b_$f�@ّ�����h����C}>��^Y"Yf�wx�B��t���\�<@NwS7<jW���S�7�J�	b�%�k��p�IpÉvНsR:��3M͎)�]J�M?�h��\k��e6G�?C����a]$�k�US����M��4�ڗ�l�M5�h���V��N�T�]kx]�Q���4��*c
�g��|<c �k�����W�J�/���/o�T�u�(��Ү,���kV�St����k��f���Z��R���#ʳ��(v�?5�\�c�X|F��z���������݇��>�on�*<�"�Ku�[����I��7t��=�[lfgf�p����p&�Z�mOƲ��T��6��1�h,8�^>��	�Ң0�i��}MG�I������̨z�$A�`�U�(P}���y�q� uH����  c�IA��M��7w�ړ�1/�v�C'g;���F�7H8 Τ�I��Ih�����VaC���-u�l_��ٝٗ�W����
�|�ƮP�j����1Lx�Һ(|Л;�I�%��k����;���}�k�j��T�ڍ8��br ��4r4}SVm����XY�3���9�P���u��^���c�tU�Ӈ�]��b9�}��V���6��ڰ��07Zҿ��T��_#�p�����>4^.n����u�w�A�"\Uov�.��h���0��>������6���@3���F��b>�(���9����-�k1�Ԫ�R�fT�eI~.�C{}����3�+5C{7g�����@����o5���0c���KM�[	ƨn�M��!�~��5Ԕ�Mh�:�<��{�M�ܐ]��k\�¯�t���ѪhoN�"z?�w�N�����T&�/^�#j�WK��j� �a��-��nf����;Q�g�9z
��n�Ãs�K݋����l2Ko.���A��z�U�)ܿ���f���*�s�Cae��L��q�^�O		���y����:��D�����|~��L+��f���@A�y�����hj�N1ڗ�X;OiX��1!g�؏T-,\�i�|�2x�S��i�6����]�:a������?5���כ�� ��!��Z~(��U���,�X�`�@�.;�w�PrR��8�k�u����o�}�
�d�P�N��X�-���f^��%�7�r���Z�¹�����C'�$C%�n��+T�Y�n� :� a3��WU�H�A4��K@Ԩ֜x�Xd�B�d��C�⟩�������m���ac,9�����m¸���-*h��^A&Ī-��fͣ����J
�,
�5��{�Q�cZ����Z�:�Oz��q����}�
�������|�WF��;TGք��m�q���FI�KS�!G[l�R����ׅ,�tn�s�ʊ�Ļ��6���)mMM���ߍ��K�ؙ�4��眓=��V��md$�ǩt�QK��?�E��2]|)�������5)��q�t�p�C­��ԡ�
��s7Z�+lH.}۩�m䏿������30(4���r���:�. %G�ם��%]�{d ���h��^�`R�TKS�5�#�9p�7�T�ϸ�IJ��!�������?'aD�h^���}*���Q(��N�*W�O�Ҷў፻�Ka�����+4��
 �ne�CG��#����� C<\5�ۏY}D
$�Xsϰ���;���T'ϑ`9,�O�TܕP��8լ:���%�E��eg��}�ϪR��Se�7�;��UIb�kk7��&��ԉ�<��U�b��z;x���N�R�3���=���L4<��K�8ǟ� MA����c��|į���ҋ3%�@ �C"��(�
F��?��6_^Y��b]i�����ƫz���^���
��>�Ԋ#TT���W���\=բD�k1�����o���g'����s�H���N)F�Ȓ���:F
(�Ui�\��]%V59���
 
I��k�+hgG,�h��M���-j�Ū^�ؠ]$|�4��{�C�tzow7H��-������	`R�:Hױ�5Uy�	��	?���B�Z�o�5��K$�_oȱ12���eQ*F���L��`�~n������й��m%c��2�nC�1s9����:@T�����s?o�bB�������{�Z��=D��@�-sFÆ���J�Hm����]�Y>D7��Q�t��d�#]��My�E)��m{�݃���s��I�V�/��Z�0�E۪l�4��?�"zv�4Ԯ�L�ܺ)�a�p �<���F�w�Sn�n����e l�wN�vPP���J��źK���&T�8�gh��C��iW�NL=���h^On��O���-��~�Q���o���j#�DX.+g���o��ɗ0���2|i{���N �!����|h:/~=�C'�`U/�U�]7�7.d��Q_`�Vگ��E��/��|�n|m�9�	�n5�FR�Q���Jm ������-+�q�Xk�J�m�#� ~j����HdHش��b"@�
'��YT=9p�\2U������yhv
��і�YXԕ��_ �z�]}ȧ�W�f8B��f�?�� ��� Mjkk������Y��}y���7�î`* bX�h�Q�$u�n���Cu�!���V�!I|(���V���{����J�$�s�x���8z@|m]]�ΰ(�fC�%t�z��z��/�޼�]�� �\�\�,]�6\��Qw�gp�?j�d��9Eg�>��YMؗ7�.��%ݱX�\��XT�%��(�/`��(wfkk�40G�9B��?�C��2�X~�\���*Ԓ/��}�]��v�a��U.�mmvG�0c�ڙ�Â-��V�<H���6aw��G�ڝǗ��.�w*�%6[{�m��"?��Gfe)��.�R8�$gx?G���|;?%e8��PT�Y[/f$%��8��޿G��Kw�F3��|������E�����PM���O�t�2H�˯]s��#1���J��P}/`PWk$(�v�G浵������j�Hf�# <�fgmo� #=���M�����\u�查���3,TF������zJ'�fV�4	d��Ɔ��?G(t*�7�n�vt*��	D��/��+<�_�{qNyr����b�1��*�Q_�[�@ɝb�c�������P#D�^�d�404O� ĴI��*~�r,��t�*v��#!G'����
�=L��mI+��g-��K�c�� ��H8Vh������Pҕ�RC�LP��fP1�%?Z�kn�~���ՅS͊� #�X�ud�(k�����[�98�,ȅ]�% u¾���� e����v��: �&��JpK$����|W<3�h%ῒ�Lp��48X`�;����	�(���a��Ԥ���hլSmN����.�h�j�Tr!06F u���<��<	͋R�_��LL�:�g@Ӣ.�Hzx�^�v)7fأc����� 7�<����|�`|i� ��̴�Ք�@��������&���;����x\�i-T,��yؙd��=p�(�^2Y��u�U7___��U^��Uk�)pZ�#�fY�ޝ|����NF}tK�a�ן�i���-���d�P U���q��������kE��

��N�pg��o�7|��N��ƕ�L�bE����D"�ɓ=w����𹅅�x��e�6F��-�>\)b|�#�#k�Q�<GhT����t�Fj�b�'�-����w��Z�?P��Bh������;��&z���+�w�Z观**^��#;��/�ɱsm�7ط�hyi�ʛ����18����
d��1�Ċ]�����)�ij�AG�>n�h��!^����s!�i�U��������M&���G6 t����g+޲q�e �R��3�kg*N3�-����9�k��������_CB7 '&^ �6����@-��T9Bٔ�lV�{<��\*����HW�]����`�t���l_��iP�ڰ=��"%U`ꢌCV,o
��՚\/u�} ���I�`"*�$T�vl�B�D����Y��#�k�}���~2����6��1��w��֏�uww������#}��q�=�ov�����m�-Kcg}����J+9e�����r�L�bT���L�����;{��uw�����n����UV~�z�Ư�=�[l��8���X�x��M�M��=��mq���ӿjg� ��@L{�/(��#B����ʽ:E�z܅hc�ĝ>@e&&���~4ٵ��	�lw��F�־B�	���tgE:����p�h۬޵e�rc3e���v�`�j�����2�<:���>���9��d���#!��Jl��&�����t�������`�3������o9��iQ�	j9��1�'�1�����"z�y�4���_Q�����{ĳ�~#�jo}Kh:�3���2677�l�� P�֐H�����qS���?���ݟ�����&��QW�~B�;�{��P7-�mycr!��71OJ�0[�u��N+����֤����`}>��O�V+K ��ȱ:>^I	�jR��t�n��r�s>�ʍoL�e�zI�^�#�䤧���3�_Ct�?}d?�@�,~N��Yh.5�1�����o�� ��wyܻ[tyI���v�0�!��-*��e�(�}���|��б��k(6�B��p�!�5���s\�gz<��h\�lܰ�j}ܗ�t<��5�#?��XcSA�a.v�:ᐲ�������:�&�ݝ+܆���������כ'h�r�B��1����hAD�	�͢��)g"¾�@:;�{x�w�̚��4o������`o���lj�[����8���Y�]y���%)h6�m6�a&��z�f7n����Y��ڞ#�%^3F�5�.��뚘�M�VJ��|�N����x�<'g�e�
�ڸ0������heuϒ�z��3c@+A����lB1��b�e�Z]s�rNs�c�������:m1cI���+��;!I}񥓢�oc�?އV_�g���1�sQfg{�����k��J1��x�X�����cSZ|�İϕ�[ǭ
��́��c��+� �[��Eu�,~������T�<��C�H��@��I�vk%���G聃���'+&�f���oj
���]�4@a����i��Ax���˖j�j������LLLjV�A�����S<���|Vw��l�b�luzp���ѣ��g)�;��K&��S�n;f�)����Ɣ��WIM�2��c�N�K!eP'$@�6v��`獵���P������#t��C��n9��>8%/�Đ��P��e}(��y��cX��뾱��}�,��Mw�ւ�U�jkE������C5��V��ho@? ��ɩfc{r�bF�c������?�RA%zhӔw��Z�M2Pu�p\`)ewWd����S�X���P-��]w g� �zM��ɃL��UT��ͤ�ٚxchtP~�66F��&3ǘ�Vm'��X��la >���8s_���q��ͅ�����Z@.Z�(ѱ�����o��ola�[k��|JLT4�~h��-�ҫ�=T�B,�9�g"ى�e�&��2f;�L`Mdl�����L+�����ݟ��+*�RN�^ˀ��d�������ag���@��@ޑ���P�
�v������$�#��tFWo�wWP�@gy��*�vTy�C��.�c4<3���ʹ�vsҁ�^�xʉT1Ћ|�ľ�؟��#"�����[D�i������=�z�����g;���H�ӷ�|�b�����+��h���1�X�ʼ�Dq�]���Ȥ?μߧ��k�	�C��&����o�Vy󹊖���!%v�����[*�U�*�P;�a S��h�Ym���w2#�����<>����w�	����$m��?�i{���E�����t$8��%y��Ob��\ll�O	N�j�.[�ݲU1%���/h�s��'r�T'�����D�]��<�>k�'?�~���꺕���Onu�&*f��$���a�?�ح[ �%�� )/))X^����Y%J}�mT���:����g��/�`p�1����)�W!*���u��CY*�c��rZ??&���8B#GLj����83t�TKKIؗ�ݫ Y-l�PIJ���!�n�UYD��8������Ą����i�}��y���0�諮�v-�Y�c����{Z�Z� T�DG1�6��O��?$�^Ze�O��k�[
�$�+$1M!v
� .A���DW�C%P 	�pHV6hqߴҴ�B�u��Y��l�8zG'73&Ʀ���ZF?E�¨UlD�rMX�r��I>��n���.��㛾c_8��=幒��fy#���])�I���T�0$������5˞�ȍ.���Š:��>p�b	D@O���H7�>�t�N0��L߳����^���u�� �cwT��G�����e��m��e}%�ɲA����09�,��o(�di��C<�ַ�s�v��=�?=\n�~�z+�~����0�G������\��\" �'m��r��@l��^
z�7�3�}�< �=d���`�,&�Ͽ�ȁ�A�qB�g>i��?�9X�{����sGGO@�k�]:։����C���CK���c&b:^7��x��B�҃�>��*�j>�%��,��ω�zh=|��`|�CB�?ڢ��w[K<W}���+.�����͌3��������ҟ�7�-�'�I��>"�=Բ{<���Pg+�1�ogGDh�S\�)9,ջ�ig{�F�
�H�h�]v�U�FA���^�<�Ψ��A�wY�����Do�@�Q������=eD����T���\�n�bB�8�����3����#q_�"@VfeA7O�}�TW���5�_l7�aqj������錇���Bem���jKLk�{6&%-`�xxx�-)Ȟ5�Af��_տ�=Z�&�{t�k|�g�=�����R�^��MF�bu��vЀ�1���ɴ�D��q���Q��Ҏ��=K����67=�Zhs �.���s'}���KG�![u�>Q��]��-���G���$H�+)x�(���f�(��)���Rn�w�)�1$���k�I�մ+\��:�>}J=�u���;n����f�� �k ��x�e� }��h�N��A"�y � ���1lw��Yj��u8���hC ��O	�i�ӵQ��&'��o7��nL�% ��rs����n#ɪYPPD��A}��� �N�:�b헀s�4���3Jw(!A�սE�\��?`��x������nx��72};���w�I���c������x5�S��޾�F���E����t���
3`zQ�����o-I(��8`lf���P�2���	��q������i����C�Y8.���Wo����s��_�2�Z���3`�<��������n�ޅz-���}]]��� �{�i���F[�@?�R��7'4Z�)���?G���g��=�ˁ'v� IA'�?a�JV"�.��c��p;������H���L�c�ss���x�Ԉ�x(������!9Lp�;�ZRR���Ϝ����s�I��f�5���{���ai�xp�i�����WJ1!��������������%�<#���AA�v�m��"�.{ػ�j�=��BE�:F�]H�����?���0�P���[d���N~���M�[������U���A?�1�$?���^�X�&A:��(Vk��0E74��'ï��.*#�����;�U�n� �j��"I��9ձ����k0ļ�&�И������)�˿tsl8�����TyR2��q1��S��y3��9�������dp��=x�\������}���#07	xE�6#����$�r�S:{��j�����;�K���P�9�1c��Ǚw.a��ۿ%u�t�(U�>���Aii���+� �UBJJ�����߱Q4:H���?��@�����IHJ�����3}���&Tp����Pu�9���7-e��h��1�}Dp/��N��"%&Vh�*y�[����ڻמcM^bLi�,��_���α��{Ȱ�#��$ov��IIe���d{;fbr�������'ؒ�xQ7�;�
{m�#���4�՛�����6���Bܵ�H�r0��/���!��vIW^�v�� g@d���e�P���" �A�r����\a�f݁2��3�	�I_@�/�߽���(��wm�����F�	@�D�:B,׀�=x���s%�у��Y��탶�l-��mHf|������j�d/x}fH��:���4�������~^��&˽BB..�~���aB\di<�L
lZݢ�-g�lы�7z��I~�g[��o�y������-�
��@��w�X0��V�^5�%�	��j0�� ��2��{���������������HD�t�޸�,��������ő��ِ��f�9fL"s&��Z[������/C��<���~l�Q�-��,�=(r�_ �媭oI��_w�t��)\D�#''g򂤤d�nw�K�1QI	��!=ՠ��{{>��c�x<�[��[�
�KU�C����/��)�;K�1�
���A\��3�+��� 6+ PMW�{zvVz)��Q���E�:�!�O�� Yq��Q7Ru�	O�&%�h6'I�[^��bKٹjSzpe����IJ�٠��鐤�r���hxxc-�/(�y�lw��B�ԩ|8�A��4�����9{DD���x
ԟ��Q_C�1C���f��15��<���ql�Qٵ'��������������0?>:��۷�P�����[����#� _�:=K'����+��6F}�+a� ��ˍ�: 髞#I4�����]!l(�:p����-�ye;L�_�¦$��f*H9��|���Sa'���δZ�_�)���de�����2eM7��x�U����5�۞��?Ѡ�.V��RKl[�ْVv���,kf��8$����y��_Y��Qʱ"�7�/N�P	�����.��1x�g���i�F=�Z�� mѯ�nzZ�fym���=z8�|&���q9"�k@q��}2����e'����=k�1��ץ͔�o]j��M4燹�1q���������:F���,Zl�wh�����R-�n���F����~v�ш	�X,X���5�z�/B{�Ą��ޣ"����\��K���� �Ꚛ��$�`�([9�]C����RGd� `�}���A�}������a�`D��F��TG�V��4�~�����Q�d	/U4z�� ����vq�u�n_�O�X�a��0&�fA����
`%�
� �A��[;Q.AC*�Kr�ah�q7�"E��=�[K"�����o��ꈲ��z�9�f�O���Z�h�"���'��;xmct�������Fi��޼��T�\22��\�k���n�����D�2Xē��e���i���:�[��-����H��"�چ�Ln�bm>���Q��y>��@�10ЀJݯ����#p��GD�P�L��O_��u�Ի�p�v��F�T
�Yx�M.�/f%k��|����\?�/���pK	�p �-�V&��j7nY\=���\"�Zs
���٪���
����B�eJC�;��0�=:�L20(;�|T���u��l�\W������a�<t�.axd.Ĵӥ�^6�������Y����ڸM�3"� �P��f�Bp�*���\����S���:���	ך�{tp=qp0	�(tƫ�Z�ʼ2<ʺ>��d l� ���%�_QQ�U9/&��vy�Ѭĸ7��{<�T)_��ۗ��S�5e��t\��s�ӌ���oY��d�����?x�Ů�y��S���%�r�Ue��>��p��`�0%O�ɍN	ڎ}ӆ�|ߤč~k�)q���?�R�9C�]�z1����'�׫z�q�l!4������l_"=��3Ր]A]��d1�n|�YVkMsn����I`��:%�mX<��$�J�t�]W��4�U�EwllL�k:�T܋H�6��9V�&۝���)����R���Fkzxx��a ����$�#q��9���@N�1c;�Ph�	�b'�Z�m�w��j�|����d)_�ܞї������pO��8� EM�$��j֚w�4���T
{����W]���~ඪ�o��\�鮚�7�:|��P|i۟v"�KP����mn�WV�7�5䏋�=='�ڵ��L#	�O����f��'��I`�t�*z�N���xn`D��P�7Ѕ#�4����H W�����K�ʪ� {"�{��
�v6}��#�|�e���ۧ㳯v��M[݋�if�ǵ6���p�����8Wk3��<D�#�޶N�k����ШZ�Y�|��3
ڙ�#�,K_m�C�����j�ҁ��̼t���{8�lvV��6�E�K��N������o/��'|��*n�\���>JY兕���dV�H�ka�;R�Ŵr�Zzc;J�J�pb��k5����`�����0��`��)�@_^����EHp"�$�x�Ʀ��v��msɌPL��/���S�8�`-���:���=d��gR
"�;��9�w�������wqP��C L�6���]<���v��I�h<m�JXƾ:?wwU���(�yOqq����2��(L�š@OV��R����n\⻎�]~��OT�q�!U�{�bT�V�(�۩\��;�Ǚ�Ha�l+��)��պ�I9<��2��O�ƞ����UJE�#$e����\���cz��m���,6���~���]t�/Pbh�[���g_ZG̙���uȌϯVYme���*��������g���^��"�B�Ԗ�x\z)�o������c�w�9{۹����ʅ.%Ͷ���ZK�*�o�W5�����M�ޛ���i��Kwy�څ���7�MB���P�%�������6Ck�����a>P¼���_���s
�]hPk�#�=�I�a�d�}�`{I��;�?����o�����h�_���Cx��<Sh��{��<�|����ⳳ���
���t
[ZW���4_��Rv��mv�)�O�e60�2%4:3AUk-�E��e���:��@��كG��[K�	��.^,L��f�n��H>?�L�Uou���O+ZJJIH���R�]��l�g�[�D!�}�"KCI�ck01J�%�c	��6���}�.W\%s��>�����rP��\�]�F1�f1��1���{�*��Q�ϛ���o6@pfB��n��:֬t���9�NGEG�WkYL���kk뤥�
��
�)?�$]���9r�Jd>��FR��-=P\3���e�~zSh�+�h��d��).!Q�������:�yI�{Y�7��`�� ��,�� +|�����u&�!"\�����5�-���_{����q�:����b8�Q[���hx���;�(���F�H�1Xz��9��s�"�����Һ�.�
Hv�������y�����`��#�D�V0h�Z ,�>��5��(K����76A��@���i���b�X�aVȢ%�N����Iw1���t�`��ݫ�,;��̻�[e�IT�� d�F����b��qɍ�K�"���]ŕUU��-KMK<���1Yw�y��y���7+���^�!�t�u�
[#7+�����G[�Ui<�6G������^�5jVἡ� K�T����1-�Õy��0$���/�l�毰C���� �b��������V��W1|mg��^���L��:^��h�/�w���,�|ͯh�N'�Q�ւN�P���=:���q��Z:Y��o���x�g�,|9���]`�������-��
y�=��ME�u�H�m��|mb��������B�K~b+26I<K��4{�ۻO1�uX�J��Ǎz�+y ���$������А@�

�u�v�. ����Vy���.�Vw�?�:+v�������ՒS��8à�\48XW�u��ߟ��$t�z�}�~ e�߿��`�𻤜xc���^��V�k�_��?ج]:ӎ1_��w/��ݲ�^��w��
>?쫝��m�c����/������=d dT2�pG�C2��s7���˗/�I�G"|b�&��G
tX��v����3Ul=�����뽏��Y���G��**��hu˭v�����|�M=R�+ ����g���/ķ�³��HW	@��E����S=�<W=9h�������p����������I�h��1�e�m���F�U*���~:�� |N��^k��0��g���]�
�w��Ƙ��=��r��Aj+s���$�	�_���y?4��6�(��%��C���4��ۚ#�ൔ�7gR�s�V����c�/�2m���󹕿o�����%�����0��36�hE�-�[��`-2,.�oWc��x#�=?r�w�Yk���΍���q��9�.7{�5����h��B��]k�Aa�����*�ߚ�u���*��|�����R6���xB��$��g�B:l�[���%���B	�S	F�z�^6��b_�G6�ȯO[���)�3R�<�����2g �hDF��?T�=v��۹x����ju�T2x4���We�{狅N�Y���q�ji!vb5+N�%�Ea	�X���ג��
;���jp������.��CϢw����^h�k�)0(�	�����x��%K���>T�s<X{��&�sސI'�d��8�/��K�z��Y=��w�}r �$zJcg�I����i��q�y!���:����5��p&��~U�ǫ�˼PMk,��x� @8�z��iJ:�J�w^9z
���Y#�����"�\��y�����h3��Μ�R����|������ʷn�je��
 ���Z�L�d6��Ae�AL4�]rnkٵ@8��`@4ud;�%pU<��Z�p�X8s���Qd�!d>�]���T�P��
r�䨟[z+����~�7k���'ૼi!1��>ۯW7��.e��d���g���y
	���Y;x;��%\Y��&� ghx���v��X��Ǫ���qY��dt!���_�<�,p!W�)  �7v~o�z����c�*��b��= Y��4�ހ*�V�A�tP��3����T/$���(꛴�膺{)a̍���[��F|SC?�'@1<��ϱp-���J�a�'V�\��Yo���y|�Y�����J���i���'�̑� �rtu���I���2���o;Mn�eGG���X�{q��牕=��J-9�e����՟������b/�L�+M���Y 0�����v��7�h��?1�W�B� �ƒ94�}|���ﰘ�!s�3Fv�#�p�E��p�� Iv巏�=\W��3K!$�p
��+{�ĉ����9+��1#2��$[)~��W�졮�Wl�E1��37S�{��l|ۖn!Z���7k�s�S�A���>��{n���ɦ�����f���L��W�ڤ�\\\&��Ft������WQ��J�fZ�9�V0V��)�]��Z3��;}?�tZ~f=jr��f:�-�+�YT\����/�g�U+YWhVS������`;����|�s�}��lVx821�f�#�",��.�/�0^,��ƣ^����;1thb'�%Z+���z�0�;��\U�p�Ω�1�F�?K�{fsss,z*"��W�y���1X��l���g\--���F��xUF�F�cU�����!�?�hQ��R��|�t�!o��諀?�ƾ��bbb�l�0�� �2��ʗ����Ɵ��������(�fWś�#�ֳ�g�;5<%�}��P׈��I�d9����7��=�bo�>Q>�����V��ipAn0�IB���+�K�-�s�vv�]m(Y$�sK�����ҹ��/�S6�ee!�:�������7N�9N��R�����NRk'��S��Y���s>�~��N�WWRr���4nsjȊ� XՏL�țl�B�s�{j�o윥����d`}����G%�x�I��Dֶ�||�����u{"ӿ���,v3ڰ���}��5$��i���������)0�C1��h�^W=�S��s�O�c��>�H���gKi�?���4Zo��kk���e�j���1���lp.�����<�)��6�o��9L�+�B�	^�S���b{�e&����Q8��Y�ɩ��]���|�1^^r����ĉIj,[n������tڜ	��<8i��-&�m���YWW#�:�ܣ��*ccc'O�Y�m�`�I��&���Q�.Kos*�jG �D�Uz�z�����!�{d}v���Xl�7n[n�b��yT��Bl��j�͢򒷗�������]�3hZ�$��o��&�C��R>�=��FaBI���H����J�)�ɘ��>�1���APr�V2���?�k{!d�{��U�ܩ %�C�÷��0��QM'B����uM��1�Y�c㤵*@��ݕN���龆�r� 0^W�?�
[ܤ[��n��RFx�c9�>��r[�
�΋6tQq���9����߾��r�ȗy���	���o���UT�N�����'t+��!�@��f�n��j�2���iii���[0e��d�|�,G� �d�8$2rǛ��~�xc;B�y�!.+�]0N�D�_Ѵ�wRCN�v;aXPW�j�4�]�u�^�}M�/?�Y��<},� �������	�X������|xP|W*炏�:��]ڰ^!ZmX����q�b���Ą�F7ʌ%������
纉�t�C�V:mSĞc�Q��Dے�ox
r����~��/{�Y
`7_�|FBJ�w��=r�]ss��A3�����n��浢�h���wJ%ee��G�N7� ��t�����Ip���wt�]���C�b�r�0h����Β�� D"q�D��Q�t@*:��ܝ��)�~����"�`Y�|΄
��֚Nn�F\޿����T�R�a3R%*�u�oy���->��1~�\���!�P�L�V��k6�'oʰA�OO����N��t
��:�nIR�<0X����kǞ$���dوf�O+�Q���(����Q�\]��DS@m�\]���K�^���%�1ƈ��jv.]	$��D��ՄL�a�R]��ع9�T[��ϒ�)�d'2�{R\q���}Лڒ�f�B�X�����_�=����&:���6iE��@�K �[!`���0J�̱��is���u�q��N�V�$u�uvuu��W���}r:��۹2	�F���.1,F���M���B��@�2� �w&�Z��8�i��������?b�Ɉ�rD�� ��ԝ�v��2�2T��������U��z�L^Ǖ��޸$��舶�>YAV=ooC�����8[c�Z��C#�������+eD�=�5����!5@�N�[�5��V����qa����e��OG'�8{�$ H80`nʞ�YdwGn�w��XB��%)ʼ��%��z�-��Fn,��Lw����"�	[A�~�h�`���O�숱�*.���ؠ���=]
����sso�u�T��!�JK������F��z�P`P�W� ��)�/r�Gi��##C�R�.aH�0�����Z���%�C�
 O�F��@���3��c�>ux��� ��p����³��p]�g���Gk3B?ѵ!�I�^ �x����3T����f%R�L	�D�Ϸ�K_�>x���� �¥$5��աX��F�j�!װ�&u]]B���<3��ܜ���)|,m���$\4ʃsJ7-1���_�82�BE�DP6���"�(�47��B]0U�q�O\��B��n.P��7�.΁�4�n��͝��K&�X��r�.�b;��&5:�FB;���94��V���eP���4?Aۊ� pI֝���pq�����������2
�����ա��dj�ND��']ܶh��y�$�ͩ#Ҏf�܄N.�G,��y�ݛ�t#��E$��Wy��嗣�=�"�(�#}����7��&%����m���b���#W9��ss�E[�{C��8��:�	=a�w�a���,���x�ދC�G"[�k��a�Ļ];t��L՞��,��tG�Q�QMw���4Ҕ:�P�fgV�5`������ǆ�ZhW�R����B����9_������vuyA��ó@>�VihT���! �u򤽝�)`�?c7*��^���#��������Y�=�,�:<��Q���r�;�����#0��	br�*�fo��˲Ȱx�5-�A��3C�}���Xc��4��j$&!?����wᠭ+�Z�:$v�ā_��220�J��F��~ȓ�V�����k ,ȗ���,B�~;4<[������ �2:��bзA��9P5�ݘb���@"��{�QTC/'ǚ�ĉ�\�M`�pE�����;���T����GNO��ӂ�WMɫ=�Wq��!�U6���}��˔�m5�V�Vx�����?�
W�ʕ���f�1%�b��sôw���j~�����;�N-��Z�ۻ�F�_�^���|U]]>�� �7�'+�1����غ���D~qII'�bT�^���{ܧ0d3C�	Z�%V���{/�o�ٳ>D�H�r�T���,elV"��>��$a����Z(\OOOKK' ��~�r)��Β�fBN��*��R��XQ��h��Ro��+�+��\:tamm!`���i�^�w�} Q�\�և�}΀��A�^��i�.��g���b�v�R�by��Y4�%�lE0�X����G�d�;����m��%?����W̑R�)�*��"�oox�������䪪���Y�U1�=�T3�X��ý��o;�A�s 갇2�2��I̍��A�
De�>,�"f��U�B�f��S���j��0�6��B�R[�1�-.t,|�?eDW:�b����U��έ�Z�z��N2��^�����{@)��}D�e͚%��W�%x� ���Xu��U)���GJ�` t�h+�K�"�zNa�W�y�@�����7Q�̯F/ '�h�,K�w�6��ro�֚m��j9�eŭW�9ݽ�ָ��Z�����T)�f�b:Pd��;���� ��P��ңV�:�'��>�y_
��H;������y���AC"��9�K��b�s}w�$�E�v���� �@�&&%�n�Ei��Z�vގ��*8�����M�������U�[��r=��<]�U��̥�얒���W�6�:���_��텂h3+���k`���rt�QLZ	�<֢�
�[{1'=��֘��?��R'&B%$�ɜ���n�O!��f���`;!�%׳zBlP!^� .�?���O���bh�s0��l�Qa<ɓ�)X{�ռ6�B�97��}�h�伛*�b���f��=j߼z%��-�Y���r}}]LD�[�=�����5gMYv����,} Q<<,o+���)�D5�MTcIi)2e8*89�����k�&�׊���Agi�ʲW���] f��W���u�-����|�;i�?�ȵ����O���%G|�76�){�VlEӒ��Eʼ:c�j'�5\�r�1�G.�&���V'7k#>�������x��[|E�d(P�o|�����A_�B�����+T����)�	Wˍ�˧��������!<� �R�i%Q���#׽!��f�w�T5O����8��l�H���}����K��:8��|]�������*y�DG��CS0arrr�ﺌ��)N��J�,U{PB|H�mf�����&E��Ez���rF�ѥ�oĵو�cf�Sb��1a:��`N���u�;��;������P�:����fBۧ���O�f%Yn�{�޿��xd�������*$�Ψ�BO�����=���T."��
�׸���LG�{�t���*3P���$�`pV]��s�]���0�˗u�B;��d�]�\(�{�6K�6s���-���5�f���kY�b�,� �ey�l��uvVK�G��:� �¿|y긹j6I�{nr��nטo�\^^^v�{W{����X��W�X�K^ޅ�
��- -�u�~N��|1�BBB����-ԧ.?��v.�+/:::�\ZZj�"D��俗|�4�#��t��X�N��)>钘��V�&�=p��:,���1E�A��7��ʉ�$4���ri	ٮ�ЮJ'�N��PHZz��NMc���P�q�v�)^9G�������R��F^B��OL�߇�"3������Q!X��j��v�눡|#!����g����4�����?C����5���/-jX��0N$=��M�{�PǀZ5�spa��|F�ِ�Ƿ���?*<�m���Y[[���~3v����*םP|�W�2נ�?c�{9=����n�X괧�)0I��������}�=ϑX;���������`Z�'�e����"�Jl�!�����<�K�X�=R�_�����Õ��|�:]\��/2��Kt&N���GG��bp��zTĸjn3l�5�����b&�¢=||
h��1$�W15W׌R�WqcR�Y#���3�>�v�L�0��`�闒�1�Mg்	��C��T�{�W*��ߟ|�d�`�Dr��Y�̸��>0�$���Ao���4M�<m �<�F�Yx`��'� %D,�R�������1�#����I�j�ֲ�+#s��f�K <�~͞#�勼N�A��04���~���j���D	ZvcZ��w�eo~>��C�K�bV&�r;Z Y�@5�ֽ ��P�盠z���z��is�Z��(ă��p�f��� g{;;5�=����&�e^ai�˸�UDH���-1H�No����*^�Q�Xx�X���ɮ�}AV�(�ޗy�\{?d�v���/�$8���z��'�ڒ�9**j&W88�Dl&��#>�2�{���VfO|̀�jhiu,ME/}�62ʇa���M�n���;ς�	@_+��@pq炓�� [Q��]R�1�U�^�NNzV��Ι��O�	3(]�N��X
h܃�n�����S�vf'���ho(����\�S}Œ����Χ�+���W\����2o���B�\�C�����܎F>�g�"G�յ��=7s0�5fB ��P�u�l(��M�XmKK�Z�F���} ��b���`�Zѳ���5�� ��_��z�%w�oq��qٕF�&;�!lQ7���ַC�V������	���K�����[�����~�ˇ����x���0R�W�3_���,����Ӆ��\�+1�#�"D�����`>���LjC$�YZ�	˧l7����$&�F{~p�MNN���r�Xzt���j6R�m��9�����T��ٓ%d��' s�n!Z���b\иw�֙39ӂ
�&�� ������e0��iii�K�Z�Kssm�Ly�]H��R��xH��y{�'��b`���na๠:����7�� �#Wc���K��B=��G!�8g�@�\F���T'=j^?�!��)��Jm�qG���5^�Qb���֣8��ք���ۜ޴�n>�`�+4"�L	+�K4�F�i<m��??��8@x�'�j���U	ߑ-�HF]���4�9x�_7I<p��Zi��\=�&==��N���};J�	��ydE��G[��i/{=`�,�o�\�{`m�E�Z�(�W����a�z����3	30�6yb�?h����]\L̬5�8�˛J� �}���� P|y`:���k�u��!>�Q�uϞ�X��G'g���$��0�C(��/��m��zw0�^���j�|L*�8�d'���2�p���?���0�U��.s\Z�=;�;�<1;77ݕF,�o6HMS�)���t˽r��C��4!�xBG.�����bE`u�(2E`)������~�G��hL��q"*�%a6VT��T��o��ך�le�$�D6±���9� 5�.���ևz;.q�Ĕ�M^��9�V ?������&/: �+��^�cvj�iMM� M��|��և�ӡ'_D����A�03�ܡ��@��H$i���3|�����@����C���~�Y:Mc�ޱ߳-����s���?�N���߷q�!QL�`��ʌB��1H	�G����!`[� �}]"���:	Eɹ���c����J`���逬Yߠ��������������q�+�G��ب�Hp��-��.W7�Be�7H�l(Ž����3��ʣ��Y�w���D�p����=#��SW{��~Te9X+�R��>+�X鬚Z$�[�++b42=+&����NWV��&�C��@�>~��~�fj�J�����7�(쟦)�?~ �F��qq ���u�=xp>g��ۯȾ���p��F��Fv���$����ɞΔ��Y)��x����щ��ݺ�R�l��g��_=+�X�:5��tV��^��а��m��(�Y- D*֚�*]�
�dW��*�*��Y=��������C�?&�D��*���-�
2
|�~��F� ]gZݷ���W��pU������;{V�6���:]/�z{��;ϲ)l���^K�fG髨��Z6f����#�����2��$i�#���1�f�܇0'�}�&�r	i�r�Ç�`���Z��D�_,�h��̙3E��Z��Yb�p�lL(�R�Уߪ7�`)��r_E
[%O��;�

[\^������ʜ��/~
؁	�P�p������[�I����]�é�1�DE���yN�� �O�
��<��H��?^v�M��uŎ(�;F졘[��fFF5��u�P?��������� ���N������?��S�G�Bq4����h�����ު�����1��JWQl�-�SQɑ�j���LKg$Οp��#$!�TH(��w�<��IX���#hi�Hr���藯ױ��cRѥ��M�������g �ݚ�_�ܽT�D����!Ӧ}���[� j�9����e8����>Xɼa��K��)d���jg�#{i�Ct���҂R��z��uz��sz���9WR�!���لh��Л�B�[�8
r;2��p���ل,qfxr,(���M ������!uZ`��h�;�i��KuEB_�D^��{�0KT���@��؞㙚����ю
qq�\�I�%&&�?�*<�W]�W?�?'"Է�*`?=]0` лp<�ւ�u%%�i
%ɖ+xl�|��''����v��7z�3%�lT	e#��*�N��l ��ӎ8~����*�;{�ZX$5<�����L��~��tu�QfJ$-	++^ ���@�J������\���`��T||���oN��8�PPKM�)� �2��	�l�WV��P���,�B8͉ͥC6����e��Vqj(�!l�/>ڂ��Zrm�+�r��ґ�����ʎ�
뽇+ݶ���!H����<G���S���0%Ƿ��ب>X�sB��t`6�e�B&tx���XOONJ-;�X��)IdJ��z�b�����*f�y��}m�O���7��ACV\��d�	�:߱5b��8 [�?_�,�ޒ�{�����2W�R�ck��V�l �D9y���I���\���L�d?M�&`Ĺ��4���JA9z��F��%�`i1�rtv6����TW��)c�ӽ����}$�%�@�k��y ș�U��� ˻���-c� 7*j�\�;V���Ԫ�
�Ð�����_6H���R��8#�"&h���9w,���>�yP`g��7��X[[��k���w;���[Y)���H�C�He�\@Nb�i�43��:��?�s�AC$����e��f�e8��È��`�Eμu����iG�і(�T��u.�����i�fck�&��fi�5��	�
�#�D�dڰ�����Z�	�����y;y�!���D�ʤP!���'����}|�������q�ҥK̓n��6]Z�I�����������=:�_H۽*%�#�����?}�]���^�5f
����uj��&F_(	�i�]r��e�צ�kK��h����#�6M��ț B��iժ2,��������-h�G��/��Z��:�A^�piX'��v��������>��Uy
kN��� Zpt�Se�F���	��u��%mٿ���m.S�2\A��������;@Ę�p��^^՜/|�*�����K�	ي��D�q}/�+{N(>��1E��-�_4(6�l:���v]�(��72*� ښ���iZ#�]��xW�dM�l��D<�fX�9ڳ�=U�/��N��3��\�ٮ���h�?�*�^�.��>rH(i��pQ�Bp���'�PS���2v|�	cK�*@V�>~DP�$�?"�&'_V�때��"ǆ�땳d8�8��>G���������8��WKHHp��= z@*z�	�b���ǎ"Lu��5��Q����,��Aw~�Zy��x]`�}�����};�㡊��$nlЉIK{�G�fU�x����|�E:��?���͛7�	I2���3H###ˢ<Ժ ���q�DɎ��˧���Q`@�~�x�1B�8������FO�s�p�^���w"�NFZ��e>VU��l4S@6�����1?�J��?��L���?�Tw�A�ς'C��
�|������{`�Y:k$R�Ģ���GV�!VwwD�������C/Oc�_���C�T	���:���{i�mN�fG�H�l]�1'ln�j��N0rM��u6�����f��1�{G^M�xIG���>!�BK(��w��o��g�N�<�����	$xp!'�F�^"o$$"r
_�Y=�������'��)�XOr�����`'�H#3~���U7&��\Q��z�'��>���ϋ�b����Y����#YԲ��i��⋠�u�u����^��������VUW=y�Ϡ8A�r����9YYV�����+�"�8���C�������yS�!���愝�לi�*f�vU�܊@�b8R��+�Y-���2A�ڟ�Xj�F����zpW�RX�����E6h��l��=�nڊT-`��|o�e��ez�/0�[�%%%�9��L���t���*���2�V������y-�IG�ť}�N�c�O�F������/��>_�|
-�_��А	�2!�22��=�	��n�=�mݍ�5(JQdU�.#����I�r�{�#�9�Σ�x~��	��,@d�ǤD��zZAN�3����������G�1ފ�2d���-���v����5r�u����MP�E~�Oډ�?
����N�#�݆������]p+%�X�,/�������TS�=M���
@p۰�q�EAU�g��&7�M^^>K����2�����_�,P��K:*T{1���Ç���)))q����5�������?=�p������	Tf?Ƚ3�_2
���hAr�QW����#�����ص����X��������Q����F`}`�<j���-������&{�XCSɚO�cT熉�y�[M�h f���Kƫ�w�� +�2����f�%�s���R�Z����(��SEqT�3A/D-��H�M1Z����r�u}�G|�"{��%u���gFbg���Gw����M�h������i�Z�n�ö��SL�?���|rz_Z�Ҳ��)hx7�Wy�`��Ƙ��##�N..�k-��Y�����/<褔+��7H�@H����=���LD���|vO�^�w�wy`f��q	��F���]Ȇ	9�w��-�rv�8�w2��,��QO��n�h��oҼd�6=Pb:D$��f��9$��$aA&L ���z��c��"����S}��.8�*-��j�-��LLV�Pl�������ޠ���<F��	�T��:uL�!Ï����g�f���V��j��,�m�7e;�i�F�333Kϙ�95�!wq9?�G��C* L� ^L�2���\���nD޹o�0r����*�@���;�{�3�:�b>�e�����ʀQ�ʨ	�޷s�w��0��d}Di� A��<E/�!�E�!p)!ezj
)Yd��>�m����q"�+����������g���9��uy�eぶ���?@VB��sz�6��L�t˚���G�]���A�L�u^�eĳT�{y�Y�^�mz���R6$�9��?N��6�|7���R6eYn�gw�NZ������M��@I�2G=�����>̌q�Z`13J����}X��S�>��mYl�6�.���ċ%�� s�����{o~��R`X���CYn��TQd��A�](6u����.{�h>*cg�=�J�{j�o��)G3W׌�o�VnRZ9���Ӽqe"�}7Mپ3�q���'���=�L�J5����;qh��o�k�|��	�������P�+�puՂ��^���6���*1�Ť�#{�����+�O�W��o��iqW�=�L%�A�y�b$��b!dupQ��v��{gԺ�.7�E��{ڝ��H6v,�Tȗ`�[����n�A��h��]�١q�j��w�pOZ?�$��g��^�[tC��a���}���69�n�������tx�DƔ����9�f�^�2|3��j��[��Q�<V��>��G(�2}��<����¢׆e�� �׍���~\��m������&w�f:w��]��{+�o߿_��{ �]��%}����S������|�V��2k�^��S���d���r�V��O�S�E�*������^iۯn����.��X}ek��=p����~j˧āCD�P��N��~ԡ�P�&��t�gO'����D[�ۯ=�hٽ�����45�O#xJ�tĊĖI�Ǐ��t��u��a��s`�5���7[�y���W������Q��Z�XWZ��Ӿx���0�!K��x�����|<=�����&��)��Yk�%r��%�q�Se�7E_}���HP=���Fߗ
��ӷEm��V�������I�b�#�y�4�Cw���o/�X�4�R*i�ׁ�;��Y��H��ȧ$Yn�9R�5Y���^J���o��3g��5�DFvh��M����15�Z�?��|�c�m�� ���soǷQMee�>[}�MBr�f�&>^o��{[G�w����t��$����ނ'11qt�ǹ�v>�۷;���)��yxZ��T�[���{v�7��J��貀�鎃fBǋ��zS�<j3�l�}W��%z4�va��/��:�7��O^y��5LȚa��^�?��|���TOXx����p��p�7�inN���$w���|ģ���4��54��1)�~���ӡ����C�^�tH1o�r~G��i��<f�r���7Y�H��gEv�E�n_lcL�ZJ�����$�n{�|n;���ܼi��%vq�#{��~78OH���q{o�/�H<�5��td�����W��_3��~���}�Q��	3&�eY�5�~�$�8�|��	��k~���J〟9��m���UEDc����W���������?�T�-a&4s)V6�#�7t�5LgЬP���&-��f���֊=)�бG-�?�<��3���Y1(��n����m������e�
�p�r��s�'��=<8�3(&33��������K�z�||�C�,�q��س�|."�R3�O��9~���QX�Ya�'<M��Oc����g�,g�;��Jw�9gn);38x�V�M�p�����~����j�)��,C3�n��1�$�3#_'6Ϭ��&��֮y)O�N���@V�՟F��b� =�~� ;�^�cn�H�:C�6(`��������� �/�B��n��((:���RC�C�Bm�Z����b&�юU&%��sñ*Ԥd�Jen�#�ee�-,�k����>�����x��sٯ��{�2������y�u^>�d�f�
�:	-���"��E�
�b���E.nn���ZCG�������u,�����lN���BB�,�?"�I���Q$�:�WI��^�ɖ��s䟉|~���w���.�
��v�w�i�w»�ˑ�1��#�N�(g��uƈ�m��	HH�x�RK�ƨܼY��}
,#���o/������g�og���A��6��v�rMH���W�Ep>�*RY~\��>��CrRz�"�a������No�J0H�hCv�Ԩ)�yY٦�an���g�޽�����fY昹�Z*˰�Z��(&���y?�y�@�:��Z |��Q�&1��|RGA�~�p����Z����'��@.����P���N���@/��b���r+=s���@��������x��]�R��x0�{,e��V���9A�Ӏ���Gz�{-1�����*��V�JZ��������?�1�6(����x��ϥy�F���/� ���;��0�fBUR'�VEaG��,�}���I��w����E4���D�_�hI�La�ȜY�"��m���u36���ϐvXŧ��4��{�b��#7�;���?�7ND�k��hjI&W���-�ѽ��[���I��	�l��K���f2x��]�y�4��K����Z_bL]��=��1��dxee�8۵0lic/�\�1�!_�^�o&ًmmO�4�l.�!�q��:,#[�����ޞ��R��(���܏�.6�c ���n�U�LJ~����œ/�ki�ڞ���Fj��Z܊k�ԗ�xrS)�jRx�36�Ѹ鷵���nxj��U�54�v�%�/��Tn�Fe��ӗ�(��\���7��ך]/Կ�`1��u�X����w�o�~|��&�����k ��ॎO��О�yp]�qK	hT�O�ߓ�\��s�2���^X𙙥\�yb�B���ƈs���G�F��E���et[c�/K�=w���1Gr}�H��>�V�����S=�p��"����	��cimt٢̽,�U���B��k�L�������a{��������"x� �*�t^$m�y�9~2*��SCj� 	ʅ�~�
G1@"��uޭ���?''�!��mL������i�������q�4�������5x���z"d�A����q��C��Y��ߍ[�T	޾����޸Al�  ��!��n�̰T�j���HLy0p���˞���u ��eއ������r��8�x�C-d��H]t�a��fc�! �/V}3g��SH�y�c>9��2��ޛ5n��}w��7�
�jHV�w\|A=���s���>W��n@����3lwo�4"�n����}��Q<��ɓ���o[;;��k&���F�[�bk������W���~=�eK��6��Na���&pvu�����F���^Ʊ�����+Jm�}m���!T�qlᮣ#G��MF����Ǻ�}?m��t^�_�A��!���Ioh�8p8Vz�ܛ^_�x�78�����h7��$�'��?A���P��>�<���-��we�%�bv�"��
�������~�i�6�z�잣�A/Gᤎ;ƾ��t��%_m��+��,��|7,w���F�ł��r�ذf������ě���1%8�SJ���]��--��#��0�)+;��y fP��tP%��oa�g����ҊG��4X�n�ڻ�����.��T��Afp���U&���W�PT�7�t*���fW�f�W��ܛgW���@8������	�,m�E�苇;ǟ?� �me̪��𫍛���I"�ˡC�����6MO\\Kmn{��������ya&%��:"{�����|��B�>	_��;0�t��Y^���L)�T&~ϣ:z���D�\��3.7,�g;~�}���mR���Ǘ��h�f74�)����o���N��P~��nΡMsҿ��b��{�,J�&c�ڄ9H�#�8��0�2#Y�?�?����y?|H��ᘻ�m-�Z�@;�IӔy����;n�ftE���4��ue���q�{�oѤ�r�\ �K��Y��@�f�P�26O޿�x��|'�	OП�]]�2\O���z\���{�贸v���H�!��u�H:��y���+@u�	_��>P�9e�O��s����/���	V�3Au���+��|D����j�<��,�O���fЭ��)���ƬE�06ߕ�t�2ɷ>Jr����v$y[J,M���.r��k��A�ϟ����ʮJ�D�k��T�P�+�Q�c����>H�U��~�@o{�FG��eT�����3/y��t�3��u>}�.�s!�����.g��۷�G��0+>ZvG�����4�����xr�Pv�p�~P �Y�o!V��q��9~e�¢C�l.5d�=���U�l��⚬j.��'�;�т٦��5 ć�K�|�y���_(1�8z��;g3�s���(�G{y����(3,V���l�&��\q�~)��6�-*�� �<ls6*M���xƳ9���z*��:��K�ΰ3Y,���_�fH��py�}����>�<��	W]�������:��F�֎0���#�i��}�^erc�f�V���m�Ko'ڮ���؂#�y�H2p��z���^9�y4�x�ax���W�%u��R�}4;{闇1]\����33�ۍ�Y�[�ۭӷn*�?�~yY�*�2zW��"Χ:�A����$Z�n�h�wc�_���y���$nA�0��ks�;�NI �C�ɦ��޽{��A� ������S I�ըy�ϻ"���d�����v����y0�$���_M|]�E	,t�n�?�afBa�t�dOT���c�c�9�t"Z:jvVW���:�2%���a��1��n���X4��9�-��i�j���;l��QTt�e��\�X�h����q1���;O�w��"4��z���!w���4��Ю3gΰ�4���b%@����h{�@�&�8�}��,9t��aө{�7����z.�eq
?�y�e���x�����h$"�5D�	���D�����cbN(�����V��!�	c/x�Tx/$�������S�XE3!BʲߦZ�":��C<�c�<�u���>���2�yi�*ZV{��F����ҡj�����)��s Mi'/Yݿ��Q�O�!�W��jI��4[!�׭�?�������W	edeoB:���HBfFd�ʖ�Yd��|#�!��:I�W���������o���ܼ���z>�������z���a�%�B >�۲����P�s� �,� !<���6�].H�/�a-���D?&���t�$'#�@��X;8���+�������������թgOk���LM��ξV��ә�t*�����ވ�~w4XY����f0�S&o�C=;WV�|�����n݂b����fnn��^�3;3��Һdh3h��8hd�U��z ��0@Ɖ��`���++Hk�]�mo�m�(��B��R�o�v�ѣ9���=�B���qh������S�z�iJ.g���}� U�J?ԣo����tV343���~L%�thH_�����f���Q����C�#uѱu�;�`0~EV���{'��~[�2ַߤi
�/�֌Y:sPZA�Ze�4���x
 8}�+�G��_Q�uw�8nke�=����/w5+���X�u�ӕ5��9V����rJ�
d��_'�re�KH���$����f� 7�bx[0�o��X�m��=_��܇Ů��o�w�z{*��X�D@u����#诤:�ܔ	z��a�NK9@R��}V�"��M"��K��'�P�_q��J��&�x)$-��U��+3W���'q�j���9��a�3�]� '����g�ɕޙq��r�{�j`c�M��Ж�`�G�NWrWj�#�i��\*!!��@s6���==�GF�o�U�&]]��L_���G�3��@%�0��Ě��b�,p���i��{�Er�l��E�R��II?�[zWS��e@�4�(6��I�8R��$�?�Er��ru(W	2������Z�}Qq�`���Q���!��7(�P�*�ŴM���ݮև�z�G�1��Ύ?	�.G��!�1�_�O,��଴>Fs�H�� �C%���ɱ��)���2��,��� ?>X���a����;��������i�N�8@��v-+s����]�����5��ۍ�Vo������~Ŝ�Jӗ/ܴ�r�q]*��˼���""�k���P����n�EtN�⡖�`��}����R���?� Ӡs�)R^�>9��C?�Һ'D"1������m�MNe^�&�A�!�����ӓH:�x����Պ�ʮG�4jQ�3M�^��+�6L\�Z��w��A�k������� ��c��}�r>>[?�ǂx�n�ä{ֺģآ���@(�l3(���1�� M�M�|������Z9+�T���1?���[l�j�Uhϡ�L�Y�h.�<��{�I��'NU(�Nr���X;���%%E0YР'����J�/Ts����Q��5���8G�I����B!���({�ʡ���%��ALq�5rC�a��T�5�&�0��A����G��"�o���ᰥ(�k�1o��GoK<�L�Fw�8�n���\�%"ϵ��ԩ����mw߁e��l�!�0�z��ήT��gB&:3D>>����oz	&�g��BCgr�\'	n�TgQUE�֧��2F5���CN�葶7��&�̖WP@���P�d%+��Dx
���z�����R�;��{��ȯ��Fړ��АL��̮G{��z/

�n����om�����C�� ��͍��d)�Q ����r���lePP T��fQ�<�v���)����n�L��p���c��&�W:	a��n�6(w���"���U�ԭ��ͼNL��Z�=����k��
�+5=;��&姅��_z�D��Fcc���,����3���47W��]��NQ���i�&���KL>��i�9��o�iOOv8ԞԠ�/x��Ƃ�`�1�c��j�i�ő�w�~`�@��Q�N[��}��z�8�v֓=Q�����
�EA�'�pm�$edex���f��H,A�Z�ܸ���s ʟ�ΐ�N��#�:�n���}�'�����JJ��[����5m}���i~���~SSww�۷��~C~�SɕX'=`�Q��ï��U{�������>�뇠�d�����re�ژ�$�&4T�2���oj:ALӥ�<����c��!i�Ew�z�%��g3��Amm׵�[�Œ�x�d�5r^ۀ_J�K	9����=���R{'�������5n�<G����+s�Lu_9��wx*�
wG^^^XT�d�;���C߀:��E��u����.��#-��3�c5x�=��}9!a����
��ָL`j�M��<%�ׯ_��tjA0�uo_nϪ��Zh���f�#�񀋋�u=�x�wM*��%z3�ޏ ,S���߬Ӭ��*�KIO/(��C�,�p�P�y⌜Q�VO��M+�vVQ��_W�}�4z=""⿁hC�@)111�B��k�!G��9���.*ڀ�	���*� U��Qg<��F�j��o���n���X�w������Q����!A�0�߿�(�[�z�=O\�p�m�!M3J�S�� P�%_F��[/gJ����r��w��hv�}xH޽�L�!����78����cܜ����K���!%
x��u@߼��Ȫ�bpp�I��c7�i[��";��J�J��p�~�qe�s���t0�]����hy�,E*��_2���'Cg�������#u�����;��Z��3�N�H���٥�9��6�$�I�2Pdsϑ�RB�QE�R�7�����b��Ĵ[���L�l׀�ba�x���u���Z����,F�\�|5w�E��ő �_0k '�%��I@nu��� H����SS�2�%��[�Y8�|J������n��q��j$~�n�/�w���j?u�1��NZ���(o�U
���ׯۜ�;j��N%''�ӑR��#<�0��f��#;f�뛍h�M��ؔnUt�lgn��,��f�?޶��j_<%�D~�>8O�[����iJ�~/Ýә�������[�3��g��3@�v���'�|�B6��hÖ)'�����������b�٠HǝN��yҟ�����,��w��x��2;ղ�{Ɩ�Tz�����/��i_����ĉ<t�UKo,�`��h0���?Y�N�0i���6p�@�M޸��BT�����뢂�<ؽ�V@,�IE���V�j9B2rrS''����+��**�>�Ds`/��'B��&b�Iy��H�
����Éd|8��$O�(�����w�.P�CQ	ķo�Z�L�K?ϯ�<�'��^��Q317gM���Qm��6��JΚC�����~h�(��H�W2�x�@�� ݫ��� '��ۤ�	�A(�$'�t��֟����9�R�x^���6H�?�00��0�!�(��?�{{�.���UU'?On�Y�Y��蘵
�ڊ1���.:��gUqG�-OQ0q��g~��C{���kQƣ�R��(v�e��*�K�Ǐ�.ɼ����)���#��e)
9v�u�I��EJL���6+�>#g��#""J��PZp�<w�*\��ל�����erP�r1ErQ�J:Y��X!饜�*��>9�UQ��M�=<�Z�̫���� ^4�D�u�e)���gdp�'�L�L�"E��f�~Sܺ|�������*�?�
'��xv�d��|ae���0�\+�Q��<�/��E{\/c,�F�WԔ�7$�E��a�I���@|k��qs0��D=������{�	"��w��l.�KSQ��Cm���K��b�v)�5\��{b��z��靝WIw���=z�?8�X~�Z�8��@��"�'/'W� g�٨H?Aֿj�o�OT6a�Pd��-�/��䱛"Lv�ަ�������]C�FC2���P�f��*R���K<r�q�7������.�m�[W ���P�O�^��>>�,Y�f�����g�I����~f��I#D�A���8\^�t��Om��`�D�Ɔ�-w~�Bssw!aa��"�o��8��%R�BB���N���G��F5�k���Y�5�=��JJ�<~e!��
p��j�a��	�Y���_�6⏸T�^DTk�0������4��/#)��cU��E����122���ʽ������Ķ���Pu�d>$�������0c�3-�P4�3A�J��䖷�׎�����^��T"۔Z�l�RR���V��yc��o���_K�K3PQ*Q�I��g�4v��u��^ryj��uF�٫=�L���F%��ؚĳ�'�#�ﮪy\\&�����Vc������o��_�������s_BZ�etTP�bָ��� Ț�M	��q��!3�)i��\y�O���d�L�\��z�ӂ@i��ݫiBr���2�&�Zװ��jkq�81 _�B��5C�㿝�#,��x�7�H�`�T���?O�ò�(�>���ϺT�4B�HE�i+Mt}�a��tI��IIo�ּ
��-=�~9��_O����`�f���z�n�߇�BC�6%���s&wL���k�NhV	s�Bx��Urr0���ZZ���6ށ1jn���&�r�8�/��{��{_?sTo�����<���#��
׳&"�Y�YyA�s���R�K���~o���h���|-	z�]T���9�>jjj�jjN4	!R�˓U_�*HBx�b�[����'��2�i��pӅ�dM8��a��;����ij	�'7�F+=�43���&����dEN�=�_���b��T R�H�g��xm�}s��=#W���P6�Mn��p�ۖɕ����Zڈ�/
C�8��y��𡰄�EA�Q�DWV��ŬF&?���͝�RX �<<|C�5��g��3(K]c2߻�+��ݎ��l��v��ݔbk�����Sl��{��鿺J(.|�o~���ޞ�-:7�1�b@K��󒷽��t<�N�j��?/,�H����i�g���q����pV0h��j��H{s��Y���uI��⫢/�ZO�C�_�D��mF<�op֞��PH�� �u�GR,@���Y_-/��,U������8!�}**�i�7���w��d�Z�����������3��753�y?�M\��c���n��}�Qׯ#�l�� ���e�G�O��/ܚ��m�iz�\K �[*x}l}q��D��5"Г�����xx`u��F�c���f�Agu9J0�f��h(��ޤD�0E����P�eQ�w�����l��oo�����0���R�mW��kN՟��%
i;)�%�쯎�#ћj��^U��#橋o ��qI������.���iC�az�����U����[���tD	9FfQ܍��j}0
{�հ�O/;�84v��adѭy�Ԑ~�,V���f��ǠN��&6}�b�@��ɤ�-|�Z��`O5x[𧪻�E`L~��FDF�����5�.O��E	b	��� A�� )�����ڜ��~��J0�ˋ�����*28<�z�3z}]��Z48V�2֒�ΝM*2"�^��i]cc�kT�G;��K���_{�Z��N��Z树^Xڷ�G>�E��R]�)k��?�U>T%�_u|$S@sae�6_���f�ձ���;��G�ѥ���BBB$zuk�CdM7 �p8M���pӀ!8Az�"at+�t�A#;;�X@'M�����5&?��Űuc��Y�<a����maL�PJ�Sa����s�r�k��'�ĎTz�'�?�<N�+VZD$��n���r����1/��dj�<sڐ��l��a��iM%w
*���a�݆�&���[�!I�8X(L-,���$����o>2�04\�ܶ���-cX��)��?��H"��o�{my�~��izU�|���k׆Xx��	e?����؋o2�.}�	TxӉ��A��0�$)�@���h�e횅�����D�"liD��hO�����3~�彈bS��߹s�$xA�2=5�MJQ�>��Ī�&C�B���W�
k�Y���ۭ�n�չ�b�}@���~1d��?����BO�}b"&���yo�,mTT��iWrZaa�И����g�f�^�l�E
;+��@:N���5��H�S�P�oݯ��#����c�t���+���,���<D���U�^nؔ|�w[1�yv����빹|@�Ǔ��� ]�p*n�:�UG-,����_{��Ɨ�.\�1G��'��g0ۓv~�74;�/��]�{�$�)�LE߫���ZC���"�#9H��7��W˻i {�d�7�5�v�w�d}�@��L�T�O��$%%��'��<h�?��-�~$��X3&�'��-����& :_k�訓�Y׸y��_�J�͕Z#w~Ʈ^BY��vui@i�X��c�t����Z�)R~R�}~p��X��P>==�@%����6L�̃��⡶�fU��S��0���h'wN/o	'C=T�}�ܔaÍi�Y�#���w�Vn[<���/���˽����V������!��6qq̏�������1�OU���Pf� <���]OIy�)�>V��k���11T(��ё\���G������m�g�n&�R'Xfh	�\[�E�Ʋa~�&m���f,a gDDD���:�@�B�1>9V�{R�������\��i��6����Z�),��9r0�&$��	͚ ��KQ��}���������,$��"�z�֙���NwD	N�qE0.*�b%��0ٚ=!�4�ޟ��qt���!���Ujj 
[�b2����7���}�#�ݜ��f�++�
�z���א-~J9��GdYY�IRmӫRR7$S���C��>����N�`����j�iT�NIi��yU8hVr;��f_�H�!���[g�R�S�QeJ�w�CP�r���v֋�n�K�
W�>�m�c]�4��iҞ�\�'�^��_����7 �f�|�=_��c2&^��-���TUUA�L��Ry����op<�j���ڜ�2E��� ru������m;;����0��#�h�	J�*�)j�i��J}�G����7�-e+��;�}��suk;�]}���� &�a��Y�-�� ������C��]5$6L�l3+�� �Δ��T/!`6�7�)pq~># D��f�]���
ٱ�##`�`T~�@[,�VLݳ"`��� ݛVy�0�ys(A(,"��%��E�Z�h��T�B�Fy�X48J�Vő�\����M1l�{1��wE�2ńU�4^��XI�9
?՟��J͹i��r��/]��&u�{����J���A��ƺ�[�0�:�i��� ���L��o⽺ T�**����L.g&����8�7�35o���
���ne��0�'G��/H��)EZ�����1�(̤��*��Bd'���%d�$@���Y���1� �[�}�E:&��hB�L~e\�8��pexE�LBa���!�0P�Q���Fk�fO��~�C��sΝ��5��?[x�}a�""�)a��@x_�����p>��)Wד�D2&��'aP�`e���r��Rr�����Prۃ+BdYr���3����ԡW��U$x�7o3�=|L k:�*��EV�0��h�У��}3��,l�į���N�?����[��"��'�:{N.�$K�0v5��@���8͇��N����^kvC����Ca^��Ҍ���%�%�7�||�ݥ=[\�����+n�������8A"p����)(Î)'S2pM/��K�7eh	�ZH���:£�2>΁`��ǝ��Ut�HG6���r����ֲ��A�"˃tt�Bt�R������V�H>×ܞ2��rRc�[^��־��7��S<�fL���a��g�O�/��v7\^ZV���R�7��J�7L,��hl1�&���,ٯ���DȡB�%7�Bj�}�Kd]���u⑾84ױ����O`�a�˻'*�f��
�y���lk������3/��Iyo1�H�QR]���$t�8�Gcd���I ���r����9�7$3��w����Xv��S�`����;*�3���w(��p��"���o"��2d@��5z!����8o��n�D��@����i�26��w�g����yWU��V�'���%��`�N�Ğ�3ɓ����E�,��ڟ��|��L){��{�%� H��f�s�-c�n��=��t�����5���k�VY�`��C9^KM�3sq�%�U�־L6٤��V�Z\��̴�u���޹g�z�n=/�?���1�긿9*�օ��:.��1	a���p)
���TW�E�b,�9xӒ��༏�ET�G1��>7X���-���0�����ݖ�8s|���Q�)�`�(���-�|�mz�EYXY�p?����A50P����\���N�#ǲ����說�������]�!'kzt�2W��9����;���ڜȈ����BQ��['N������Ρ(����&�'���$k@� :��rP��Ʀ@!���s�I�JP�i~}�H3_D�ךۯ6�P���SE��J&X�[L��z~U,�)`	Tb����&�L�̀	m3�,ņв]jņA�Q����f���<fܯ4��V�Ūh��*'L��TL�k>7[���ih�w2E���j�$��6Y�	�7v,���p�{�����_uuQZaM�k�!��SNFq
<�w�=G,z��B���7ksČ������rmꇐ����Z��?	b��% �Pd=es�G�K����������H�U6�R��,\s5�
�Mlө��/S��/��lū,��a(���TK�*�Qة�*S��]��)xWR���6O���>8���J_���fY�Nv��f�cӬ*��M�s�K��iO���щ��x��0G+K	��@�j[ �.�U����ﶴ.�����ih#q��O��"���ϻ����s{�G�w��B��1�9����O9��%������>��Bl��8�M�[�������f�?�wo�Bp��_n�>�fh�.�kH��KD+(���W�sNUM�|7h� �8Y���*�U���R��WB<�m$Y���q�������?9��ҲxC���8�@���j�ӑ��A"?�1%���9NEjo�x�2��a$�7";��mٲ.$b�XH+ҹ��3aq���H�sT�iݓ�D���h����l	p�m�,����^QY������8�T�+�2T���������� �[�8#�<�g}B��#�h�����
�����}]�����Z����+Sɩ{� F&'i�v�]R��?�U���������Г�� ΰ�:Q�|��gqq�,ll�B]���О�ɬ�����Y��{6m�KNNn���7;H���ӈsa�"�X�X�8[W��\%�QV�$�x�c�r� ͅ<��U�k��'�D�6�o����!��s������A�<�Pup�(.ʹ��L���P��͏SDP�Z��К�}�I�#�O�s��_�z�O�|��e�e�VI$�{}�.�<�2�I�p<����{ך[
K	��W��`���L�������(eS���qZW?Q�GZ��%0d�F_W|��/ ���J���/��fWa.��뾱r�kt���ĺ'�R�S�|�VW�P�c�e?��7+��IY���,�LJ.����PE��!�~`P˽�������P���n^E>��bᑑ�R>����ݍϑ�'k�!��4;+�U3�/�	,;1aJp�y$?p٩��+��gv.:���� |1;�i�y(O�I���#������|-�XH/6�H����(�y���|^y��J���ᚡ�����N��Յ/.��A$�#��W�)	�vtI�yC� W�f�jО\]'	n��{�=���[����p��ӭ#5�Tћ��ڨ78F)��f���w�&�(2��4�^sO�ܟq�w�`��i���5�Gv�H��4��TWW��(˧�໕�*�iB����>Mf	��F��o�dJ��9����;Z��/��d��Xk�6#��/,�K��!���w�1E��fQ�dA#&�#Z)�����ץ�Ɇ�NJ�~�8�4����\L�{�����4 <2�;��F	�p����җ���qy�G�|\U5J��ob��h��%
��d``xn�ğx��M��9@!�Ӟ�W񺁠8q����@MY���kj��~��{|���aw�͊�Kv�s���2�/��P~5y�:����2�'�8n<�#|E��#�����󏍇��T�a]+#օ��\��[�z��K�ꍳ�ڤ[��f�ÌoX��;���$�U�?�9��V��yu�G��}��u(r�R���{>�2�ݿS#���=��4)g�3�̦�a�=%�������[R�o_��okm�t�D@������ͦ�4�k��榦��2u1�*4���%����_��2�4�����~{$��B�;?(D#��i]��\L��������㓧c
~Q�x�U����"��nP���9;*�~�Q��N��!�����V��ˤ,�։���Ndiha�/��~�Q.��G�X_{��Rbv��"�뗘�7e�>s4&'�� 5	��%>74�"c��n��y��K<n�]^�k����\�еk��X��V��%p�H�Pu���s�L��ڻ\�W��6S��+F��MSH#����e�j.%Y���%R��dr/��_����
��Q[W]�˳��YH�6!���$,	���-Rl&?�g�wԁ:�WGQ32Z�{����w�[����ǀ_�Uv�33��d�ls�j�
_��_)�b��.)�K��]؞ק��9Ԩ�1y����f3]}}d�LD��S�֛���;9�+e��\}�"��tpp���'Z�t<��`w�#�tz����|�bz�h�v��A��%8���c0�]	)�r6�u�`hy���T�A��pJ�� �|ᙯ�Ț\����aIXq����	�↛;~�ylс�^�ecg7uw�mͣ��
<yG���5�h3Ҡ�S.��&&&�01���a�N]�����J�{��=�B�0.���U���-?����meo��%6�7'+Y�Vn��Z�Ą~B�y�Ӻ���ǯcbR*�~zzv�D�T������|����  ({~'8�W"U�{��q �BX/ �)ϭwȮD���(���7jjj%ee#;�=n@�X�渋Qu�r�HI�!��W��ʨq��X��gώ)t�
Z��F�W&��^�t����V���� �S�Xs���%�*p�n�%Oת�Ɖ�(�j&R��0o00/:h�k���;�o+�!�V]�ٌ��,��=$Ğ'���E޴��P����+�����3U�;�L����)���4��PUV�ΙB����&��G6ҽ�
���F�bH�F����W�������D��_������Y&�=�-�@D�YkU�F����c-ܡ���x0��r��b;��#��}Vw<�(�`� ٶR�J�X��������Urr�k^~��i�)v�H�<k�Dl��O{jM���U#�~�:U�������m�����d����w���,�?�"�(��+6碨
:�!���~s��b�����I�����Y\k�����Β��RR�����Ƴq�+����^2f+-��{�URۃ+W��9eՀ���#�h�V"�B�ND���IY��;=�	GB�����aqQ�f����E�~ݳ��J���R]Bc�d��\(��~`�Zf�L[��N����^`���ž�a�\�+[�ω&c����@ϟ?/��跢���p�U�V�d���2W��m�Bs=��.���2�(�z50?�<�桴1o\KK���G	t��S�1�+f���z��-�����C�%##^�d�ݒ����� d�ܮ��L�H������X!��)��:��i��{UZ940z��KetO��pŀm�\u]��6n�Qo��Y�����'V�;P��[+.h��\�eVƖ�5��$X��:9��9��o��wٲ0�T�Q���*b������ܯ����N����IG@.�����<0�̭Bdo@x�sʾ�fB�][����L�X��t���>�6I�Ut+�����5U�!���~��[�`�_|��AKE�r�� Pm�U�᭣
�G����o��ZÔ����OB+�J����M"Yt�l��%w�T�A$������LD�f���A�)��gl��)�*<������RʕLL^�?5�	��t�MRjj$���(�P������N�:��201�7M���4]�e�K�Zj�� �R��tc�->��<S��LyK���I����,H]���"�U���v��N��T�Q���4u8��N(���5���y㽟�Bn���d�x�����M���y�����6�>�~��`E�������ӌp�	�������>�:M���_���i\Z�b`O�9]ӽ��3�~�A�9R��W<}>x��Lक़�4�݀`��>2G��h�JY��i<><�`Y/>{��ԓ�I:6�=�0�����G:Y{&��9�|ؿ��A�wK�L�����{7��zV�uN����K�ld��7�9kw����#p��!�4���ء�%OO��GN�/Zq�j����a�1�B������z�� =������{_C�����4�>�2�����AI�Y\|�ך����+��W�[���O�[0^V�98R��52e��m�ኩ���`0�!�u��,�����Y%Ţ��dM[�G�k�G������F���s�t�{�&!�J�g~�FBJ
o�/kЖ|�`aUj�ˍ��������p�����^��?�֢�˹;������@a��w�o���0��K�d�t��G��D%J#_*¼Xҁ��e�Z��*wzg���sK�Z�+:KC����:}���c��C��8�h��|-j`;Wz�R���])$$'�2���LS\�ڭ��ëN�J�WY��3IC���+�{o��Vfse&ɉ2ٸ�G� s?檃��s�i%���)�>��:����/�{k�$99YHE�Q�0<����|09{�R6���9��s|#�-�t���DT�����Y�X2��mB8E� ^PL��?#x�rq�2X����c��*�O�Zy�۫1�$�����ln�9=?���2KG���%��I�G-E1�����m�� �X����t��Nw��T�kkٿ4	�����
���`̬f��|�=q"H��%
$@�-4Kُ�9g;�wt f��S���2m��[:@���7E�a�3�;����&W~�.Z��ҋ�x������ Y���_� ��>5#I_���o ��x�9
�_&�/���mtO�2�L �	*w��U5jT�%؋�J�b)��(s�8}=���}M͵���Y$:KWVN����^Q�A^��g� �0�(��7�`"/'ssW>O���e������B��Z^�>�|���,3ٛ�Ib�++`q�.E�	����v�<���9Y���E��9'@G
7Mؘ@�	�	���}�;/�@5�����>��չ��L�֔�\0<�"NB^�PMqT.�����o�[B���U22;��Vp龍v�B=�.�;N��,,T�l6]H���\�,���%w�������9}�4�;$��K_�&q�x�D9VRQfuM���[0�Ohl��+�11���
G9޸����JJ���/䢻�9]��$�y�(CK���~�.�P�?-F~u
�;5U-1ND[N�1�Ի���15�_B*�$E��A�W9Of}+�[�LML��x�IoGEG#ۊIy���ee�	֛n�]�J�#l>x�#l�2����e�����j�N5#�b�}�P 1`����D�
�<Ea)	���d)�
�$/9¸x=��n�?v��[q6��jlu����
Nzu��-������&I-~W2��[��((Ƹ3u���J30א�U��>wf�KR�9����9�0�(��ԕ+�$�M	s*�O?~�fv=�jU�(����E�$]c�[(:�'�\�F�οS��T�2���<}u
-�R��[C�=u������㩚�A��wO�޿�������R0�]�kdg�?&|kD��K |�3�z����ۨ��~��m� ��(���
˼���F�ˉ�g�����i�}�����S�
ى�"Y�ˣ��ߓ?�Df�����z;�rUG�.0�����jt�?X:�Lڭq��˝����b�*��C�Ρ��NG܄�iP���=�����>��k�֐�ly ?�|����L�+�~;T�lj5f�o��Ö|�X_b����q�����iU�}W��d`����upW��p�몴�Zj��-�~�ڊ�7��-Av�~�zE�b/$K�F�V�����ΐ��^*�'�Tdv+���p��ޘ��N@�=o..d�0 �+{d���}������DG΍���ͭ�uT
&V&o�Ӆ���^�P�&�����P{���Z݋�9����uv^ս_�W�p}a�`��������b̋c���^��ddff&�h�0�0��ں���m�J�\O
b^�\JBf�"*)),��&�I9��T�����v#4M+�� ����,��M���1�ŗUh���+Mi7y��vL�́:U�K
P�+����a����j��D�tiְq�J!d�{҉�Z����uk��BH�ޛ�p����hv�V�����.����!�^s1��#j�wpITelJ����|�L@&?8�2����C~ Vk�Ό;U����;��HzR�=�Pҭ�}�w�:j}]�'��l�0j(H�11C	�j�	Pqkj�J����{�3�'?ٻ�����˴�y���徛�k��%��{�%���_���P��m��M������n�3N�N!���C�.=�����q_�T���O˃i6�p��s?~;]�{�R�������',N�~?ZC�9ȴ��Lx������{9i�Du��K\��.HM~�a0�OF葵�[2���0�f�k_�� ��F�MKq[HX�X�B�fI���ْ�� �0R���Ȏ#��#��O;�ږ'�������_ݝ�ZF��ji7��L�,�?�������t��*��>opӳ�fKl�I�)��f�����^EX��	d��NPu��f�
�5?'@�~���'8
s�,E�ݠ�[k�E���z���S/����z��s��pRB����i׽����߃6Y��!���C/;Z_��%�X6�OQ��OQE�wģ8�"U�I�t���f�:|��g������g$�n�AY(}���@�P��m�ߢg&���Z�-:y2���aۃ�yYC��3lR�޿���V_?��^�r�c6�2�G����H{G_Z���D,q�UXb���'��[�^����hkʨr��(kk[�B�+$�Z��Ϟ2���ݒw�Hc/���]�M��l��p��$�=kGj�Uy:.��i������V5`?��ӀT3+	1+yz7>Cnf���J�uE����؃��֡�v�J����;�<_�}�-���kk���-�\��<	;��Ɓ]Oפ��x���}G��.OI82�D�{�I�#8Ů�k�Y �U�����R5�g���-�w,��0!'
==.#����	_�妺֨�GTU=	��m�8�l�?l0�b�C����g���.�����|*����J0�l�`")�}%i��ݽh�+&e��"!2��&!2��c�}�ID"*�&uz[�;c�K%��ȋ�VSI��5�P>���Eޞz�ڸ���ޱS/x���[�+���x�ض7|���X�I2uEfaĆk������raaa��9��7{�P����<0�{�sB�6�ԕZ�ʣ��
;s���i4����݀O��%`�~�Ђ�D�L�[�X����:��1�e�K��Ho�
��@!�zټ͊�σ�L�)�O|��:�o��;z{?1$��� ���QH�gĳnF��Ֆ����z�1��)������\��v�C3�Q�ìˉT
���T���z���Q�Z]��^����K��^�QB�q����v\1v��|�q0����%+#W���2�ӑ�M�'�!o<��XH�c�; @�?�"�,jbcC�l�q�=/��%o�v��R�Z[S.��:i�I<�\8�st�>�f�+6��'uk�~�"�7�d����WiR`�9
Uq�n'FK`k�uL*�-��[4=�9z�����iik ��p��w��DT�,.|Xoȳ�VVQ1�j0�LmY\;}R���Jp���	��̈t����\�]�B� �o���۔��Xe��/3�Zn�\�������~{
���gq�6]�u9�$�3������7���8� �7*���Iz������Wii%C���xh��녪PRR�:�b���<��",$Ͻ��c��࿷�֒��]�)v�M���L�M�>kv�����[k��K`�<���l.�<��q@�$������%c����yQUn�&�9���?
c����hK��?z9�@#���:���Y��[��2쳰M"��89�4���5���	@��ĘӞ�.�&K���n��.�R����݀V��F�޵B���Z+��WR�T{�n5'���H�n����ӂ�'
*]&��o:�1�4D��ol�ܓ_����\X�
؂<*yK�+sy0D�P���hf|؎΋]υ�O"������E��4
�G�M�`�"o��4~�<m�𻶥��&c<rԞ���	yx1cSΤs�^?�M� N�cҾR�%��&�bh�!��|+�W%o��Ċ�A�B���`"\��;#��g��_`0���Y��:JJWؒ_z3���J�b�9+�}몭\s��44q�<�<����9`�f��d��������h�꓁z_3����q ��A� `��-�x�NZ� ���sH�<���C�=���A��tc��M��ֱ�������Aϖ���Ť�]�jЂ�<cT\lo���勦��(�{���vv�Q��,߾��+ѵ}|y�(,��̌��g��=p����p,t �O����dv�k�r�Så��{���ϔөx��3��$��80�.�]c�
�IU���\�� �wrЦ2o \��ݳ�h�۱<�U��_�.CU{�tN�eTu�}kwwiv�>��=�6�}CB������!�w���O���_gP���$�V�9v��iy��g% �����Y��Q�MNղ�Sh�ƽ=)���;Pj�����#�n��ɴ��e�'�=�'j�����iVV��s�O9H%Sӭ�G�
zN�2E�a͍��n�n/,����BN§`�j�v�:R�P��q�^`�cBޮxH�JJz6�`�����U��k}QA~D^[%(���Ţ�QNCe-)�e��,������)3Z�4A���)�����ހ�Q9V�:W��"�}��zj�>�6G��;X3ť���W����)�ݣ�r�"��C� z����>��L�nIC"��r��du�{�H]��+>�M1v|�sL�W�4�z;]��:?���Y\F�z��ߩ��Q�o�x�{ҵ��"9�����'B>`����H� �/7D��丼��$pGHf����k��CZ'/*���s��[�>{r)>�l�u/���c	�~��h�
���<싽�| ��+�48#y��1����H�S��d������9��Vie)�;d��~C|�Io3����KQ�?{&ո���
XwS:��L�<_O6��f�%5��}���e�\ͮO����������t�������������s��iO�M;�M9AQ��m���V<ݟ�+.	~a�b˳��Թ��ͺ��ע~�T�No�p�bzv�	s��?l�9/���Ae�d���\J�����Ks�����'�i�ro 4$d�+8�Ril�6@�6ޜx{�Kct��JQ2]"vۥI��罗'ʡ�JJz����C@os|u���G2�c��� O�V�8�(��O��,�?��������i�8��&��RP�z�r�|���N�좲�Z�����I��w�[���2���������MrO����n�u�i6}��Q:7��)�Rf�$�(�������f��B����@�?n�A̩�h$�՝u��� ��D�?G{���7c�^0�t9�{Pf�$����(ɱ�ߣ`}G��}A#���NU{}��ma���;W�6����&j�O:��t��">#�^$才�Ç����� �����U���{K���-Bv�^�++�쑄�����G2��d����������x����]�z��y��|����z�^��~�n�z��|�&�n�	3t���1�5X
F��:�ʊU��Z]w㤉��ׁ7:8�A�l��Ħ)s���B|= *���(S�)5L��K�{�j.�ӏ������Y>3�s���؛JcE-����~Qo3wy���@`4�8w�V�n��ߵ�ˠ)�7�����)�-��,��7���УZ�0�P��]fH�Z��ĤOGB�㍍����Juuu@�H������^���?����1�:����������{�P l���C��21���mDZ4�R2�c�T_���r'U:w���|nre��r�*Z�O��:N�Q��.�R\�R*��"�á����l"��?ɾѴkl�{xE?>YN�̌̑,Hs�1��Y�W��uz�6���I̿C�wR�:"��h���v�.�Y�`��Ĥ�l�- S�( �x3�g~�L�#��:�����Z8c�b����'�C�����%�p� �TEm���~�O��X
��@
 �ڥ��4L�-y����g R�t��K`�9`�%ec�E��\�gh���sd�]� ��V��ɯ����.X� ��9�����]=��5D�>����t]���߱��.����|�-�睹����MMW��j'bq�s��Vō=$�H���2���=�.���s=�<H�wmep��������eD2DB��� ��,�h�/��/���|��f8L ��i?����sp(G���+d���E�����
���D�>o��������#�/�p��P�o�0?⣩���e�����ѝ�w��Kγ]3���hXb��뗙�Tʿ��XY�nk��@�NG�+)MA��fhFWhjd��"^��T���ى�i���@'H>��L-�Ő�{$,(�����Y�k��+(��������9Z>}zeii���
:	�A�������!pQ11@�y���vx]U�NI�.�w�ir̇��tO�n�hVd����҈T��֥����ۇ�[��q֓_Cer�2�8ȗ���J:��t***�?�5)���A�%�s���γ�h5�11�6����2�p��g� �ˠ����a��틍-1Ƌ�-��U]���D�n`�y�2��e���q�I�����������e͑)�H�ȆD(��َh�Y¶����Z�^�׋p�Ċr`T��_&LuV<�./���sJ��1E�����D��(��`�s�amړE�,4L�8S�8���r����#��@Ɖ,L��̸?��n� �����IZ�?;H����t��N�#*�N�>��\ %���aEjP��ѷ�m;��R~2J[��V(a��jE�6���L��3ۊN�À��],E�]�T?���?���z�M��t���Uw���j����ը����Ǉ:>���f���=V��5:Jm+�-B׊���/��)o���E��郗%�T��t
\�� $�z�#*��s����bO���u㖇��6��_3�r̦VaajC��"V|����q�	uuw��,r��31=�K�\k��H�s&7���	����EsQ����0���N	:��
�.H�r�X�께p��UņO��y��~��j� ��T�FJ�������X�k�[���Wę�ݼ/��������oO�Ggq��8�L��1��s�����Z��>C������0��[����i�������HA@�R���?�`��Բ��/ǆ���H1 �Y}_}o���(��G	JK���dJ�@�0�����C>��>0,����VP`����'7����n�<G�"x�7u�ʣ�.y`��|p/�����S� &��vw8�OGsdg��
vyXuC�K96m�ޅ{%(}4�;V���9 H���)�#�@Pҡ|���P��������{h셜TF���9���/����{�1�Dl�g>O��v��>'�}޳`�H)�{K�`@��Sr@8_�۷o�B���A譭�wX/񫫠3 ���O���X?���gO/�_��G��.c0U�!�:�=��tm��S�y�<g���3��\��@:�&*hiYH-y�"��뜡����K2�;O�	5���!|24� G�邎�,x��0e�����������]��܈9�OI�Y�_{<=b2[�z�}. 	�'Ř(�y�����@�2&Vf��F?w"��g}��#Ihxy�7Q���U���|����z��]��V���;�#-}������y
�����ҝ����/��(��Y��j�@�ͳC�&�].M��EеB
wSJ�,�ISFF^i*0?T`�ghs����t���pqO�0��!k��o�j�X�8��|�����Wn �l����C���F����'�9L�=>�À�y5��~�%Z���j��rmn��?�9u�T飒����d�>(~55QA23���f�eq�f����c�HY���[�]���o`�cx�[�������x�sV����:�Toan����^���(D��	kc��I�+�i�
:���e��S}��a�߾���Qκ�du�r$bS�w�CUaӽ�^��j ��o�;�&s�ҦL�E��\n]'������k;�&��mqqq��|�f���Κ�׮�KI9��8I�'�Y�?<�h�:����*����W ��mYY�!oj�� ?+�ٷ���)S4ظ���e@@�YR��@:r��1� qdnsI����%G-�����TW�vxz�*N�H���2!/��e�C9*��n�̨���\��o_��dk��L���)���ze+�ƭ���Έm��s������?�����(���L��O�?~�n�	{�
et �Q6���޴��9/���'���B��A��y�noo���B��LrJ;�@��!�����؆�M�����	�{6����D��G
�Ϸ����J�k'�sMinj
��/�Л+)�N\l���!�"����<���!7)fcCX����,@����S��1%7~��↳G(X�_��U���f[���²�.8b�Y���@.i�\[4܀=������2){��>&��Z��EEٮ9��s���p��s��n�a��-�dR��ӿ����gv�˟��E���Y$��r�L���|}�**�D���7&4�u��^��Qʊs�����6���_�;��.i�\�$�ɕ�_��NOO�9a��@���M	ـqS�h���V�89��H�W��=������u�J[�/��G��Xn�?Y��g�X���_�[xV)�}@􆷵�!|������!�:l�6(=�Ur�O=�x�N(+�@}
�6N�am���3Y%=K�s�熬J�f������F(C��Kե�L5`���Y�V�=!w�	�����ɻQ��_��?�Q0y�����4�W�ݸ�z�\k�Kd7�E�wnu���8�{e)�#KJn�]),����;B���:��s�HQN1*丢�b��*Љ�/��&�&m��7�"'�j����!�b��߁�����w�o�鲇ؕ�%K�bOU�ggy �1�=rx^�Z	���f+������.�-�"���m��w��BC[��=E

0k�캟����}�����,8j��-l0�G��5��Y��h�	��)-�P���bL�ܹ��w���bw������"G��1�8=�����)�Db��{��
(�ܘ��g�2��+qW��h���� ^�ҒΛޅ"Y��$��Ç�iԽ�ː���TR�%WWW��Z���Z�FG_� Q�,�!\�9��OZ�x���Z��v4.���f�y5z����{d>Ϲz�%�X�Cك�kq#)q�!gu�m	B:p�l���x���4P��-�ꅚ=%�xע���OꌡD@�#E	�Qv�O��������x��.����l���ɉ��f~��D3���P�j똚�jk�l�*9y�b��<oj��Ѓ���Ҭ�g)S���! �0�}�h&�����F|�O��z~���<��sl[KGx���5F��Up�+�5�7o��¨U��Ռ���@]X�<5/`�8)r<�7�B��|��.��'�:?Y�}�u:�%;�� ���@��O�~�6�K�!��J�i�D*7��t��uZ��˅
?�'�}�ś	TT�l\Vpێ�2L�	�7�4ܜ��n���;���ə�z��I1�4���H<h��4�XQ�xQ&�W�T�����KP�G������ӱ�F�}ij�E/l?�XU���$
�LYF~4+9"�m����ש�C���a'��0���0�e,��R�@�4�`)@ɾ�E�d���'9�|�h0��������øn��:P�����5���%;/�oM=ܽ�\��^�Z���	ʼ��pq�2�{�;?o������d-䟋B����%qiX-&�D�; �͓C��=�$��xr�}^j�5&ff�-�^?�����)��Y��r�T|P�Ql��O�K�(�ݿ��'��Н�V6�μB<�n���W"r���=VA�yC/x��W���a���9/�)+k����oғ��	j�
y�	���Ŷ��^L��(��`���o��6��rx#-Sje;�(���/4�6���\������I�tOL����HJ>il���D��AN��QEy�\\\�R����:���C@ְ3��U�1�8�3���&U#��S"�]��<ćG�Ľͺ�Q[88�B�s�ѱ���j+v�{g	2���m�uHȥ<�o��{{�Z�e��I�$ht~�wA�]��z"m>u���1�$�rݸ�����Ѕ�̡�;ZP<L̄������f㈿������_Q9�x叕��]�h	��Э #����o��gM�>��S�#-}�8���:�{su�P�К��ܸ�Ljo��8*Zu֫��g��1RN�yv�|�ghx�B�^oz�w�{2���i��%s����*=�����\���c��<(a �A�!��=��/���x�0yP���fi�(#S,R~)�	����{��A�c{9���xP�/xe%���A6���>f���%~��I�U�K+��M�J:�!�I�����z�LHXCO�/Z�9�V}%Y����������}y�.�cඉ��oK��G;w9��y�fd����\LA�k%ā|!**��4:kx�̄;EE�A�ϷI�#�Y�� �i	}_�v#VTx����g��HZ`�@���G����J��ϟa�9 �̮a��z�����W������h��M~*�S=/��	5�<y�2Ug�N�,�C��vB�5���w��(��*�U0|�pʯ������w�
>�ss����N-���hW��[{�sp|�����6@�d�tKg��E{��Ւ#^���<�m������{�A;;_QU��4�$ޜ����aw�:&��z�êo��$*�E���_��L�����HP���&�!ߑ!��Z�*��aO\�ґe��k�"��'�G��\~���^���G#yR�x�ī�3�8��S�Hz��R�a��Bj�H�O��E��~�T�K�Ջ���>h I���B����9�w(��x��'������E�؝�
���:)t���	�s���D�+?��f��IJ��cl��V�� �^\ģ��V���ua�����_T=�
��l�Ƌ���0�|.ךxv&�Ńx���r����t���P'����&t�8�������'� ��)q_���KA�'��	�̄���D��P&��1�����Y.01�$� ����X�T��@�OZ���@�ƂB^��	��B�99n�Ԏ�2��hDs��A5����,,����~w���-$�� �蠂�w��K��.x��?����=E��wx8��TTJ�xW@R���5�l[KT��ݦº�����F^��Ew"�oP����^T��L���?;���/��q�ܛ����B^&W�T�IO!�uś�%��4z~R�@��
��l���Y����<VHA�u���_�{��YJ\v��EɦS��TgζbW���:Y����*j�`�����nH�R��Ֆ߸K�ᠽ(ݧ�����Hԩ�m�{t$��m��������I�-�?wvh�%|2���Q'�ez����	��4�d�֯��p	0.P[�c�XR��Pyue,Ql�vC3Eo_JhB�j*�{���s&��G�O�~9��w�`6��UVH��a��<w���G>F����:E���Vx���FY�03��R�֖p�^���b������)7�nF���G�k���#��#�e:;7A�0��n�ʌ�+�������K�Mh������6KJ�&W��Ս��@�R}�̮ޘ�|��8[��m�QW�;��/�7P�j�R��1�-���t���'�7,ͷ��PlZ�Џ)r��~�>ˊ.����/2ά�M	7ZA�+W�\�E����=��0ZͮRSR��R։"F�JbM��.\�"q���4�s=we�z�&�����q�řĦ��y~���aG�*��8h��٩�oG#c��7u��?�(}����f�ۺ''� �$U�v��&����yNr{D�!NN?ad�?�Q��CT��������φ<w[[�n/h��@]t�7W������[^�T&���1C�t(�t��n��w�束�N�p=���d�4��iK�Á�����Ev��]@�鹽nA�gٚ�GLb�6�4[��9��&~��u}��p%^-�����N�q	�X����`e�V#������o���W`��ga�����[��geq���<4��\d��	Vnn���6��wh�`�`�y�� ��*����B��,=��,�r4���r���b����s��>��XҋI�Ƨ��G�� ��x#��9մ��+��h�N,DCHo�wB�n���4�-���������=yش��qh�;d�o$I���c�x��t�dE����j���E�:��TA��^ ��+���-O by�RI:F���a�Z�|�:�;�4����)ǯ�z�����p�q����PQE61�6y5�b0������Ǹ�:낤�ʭ�,\�8����Q'!�8�K�l�
h>��N��F��8��vu�<�quv������.G���Ø]��Գ�'
G�Eu ���DD'�o�>:�y|�ʚ�g_]S�����Vi���VWwwMuuDM͝o��5��fA�T�뤯�()��/н9��C��y2�G�����h�D�p�e�?0+�H��dH� ��q���P��0����G󾚽���wY�x/�s��Wز�ڗ���;�^���m�Y *o_>`��>����0�Ɨ���汍&���i�ts�����<�
����\t��*{>鵴�G�Y"���������z�k�>� ��8ƫ~�q��x�B�U�:��[�K��"{��MZfO��w�݋<<�
��Q��Qо��uLO���c�Ѫ@�;���s�I���+2��ױ``!��(�/4�8�R .֦�x�$�����b���̜��P���Vl����i�j[*������EZ�55
�H���r��^�ٻ��载A�T�Y��Q�zE3�m����!�3��o"���2��2@C�@R�K?��B�� r�_�;�����H;;j�ܭOn�:�_���!�G::��\_�20�ii�Q����b����`z�ID��&��g�	^��\4�ZOC�wG&�$O�5 ����� ��$B��a���m"hl�r�jn��T�����?� p��ws�AyGG6�Jd8U�x�Q�|q����XQ1�1*Yl����s�.p[�����Z�8�`x�ocZ��J�f�f�}���h:65�e(�	}���Tͺ�N��=��e�R����bȚ�~�i����Qi��ʗ��
�����+�́%��d]óm@"����H���rw���Iq	�2Y+��K��
EYRF��{5~�^�+��{�s���j�x���;��"�bG�X\%���%g�Z���h�za;�>������+����F�
]2Ck��OשB�����d�၀шB�8�!0,��B}�]����.������ʇ�C[^��[�_��(���ߖ9�*�-EC��Q++�H��<'�WQ�*%����
t��(�?�:	�*:9�`u"s�\K"�kqQ�1��9���}�]��ZKׂ��d��ß�y�������먃o�_Zg*]P V�v�gz�u�<���w���yh���2a�G��<Y}���lt��Z�x�~��*�>̇A����:�{l�AJ���61��{l�?x{��$�Fz�U@����ʧ$��۬eͫ1���4,Nva׆ �v�5h;=&��tИY[�c�t��@݊���T��ɓ,J^k_\P&��Z��׬���q?�&���%���?�#%��	͝L֣Ňn����\wuo�5�E]U"���ż9��LIDe�>���~�)M2Whk��%@X� ye���;Z!��N(�2�\�����p�{#�%�0WUt�̌Q)�B�dk�X���[�Fme�H�����A:��?��J�q��� $Oͯa3��l��ͽ~N��������Vw�t�1�r~)�����b�N|��cc�Z..�:��4x�0��蹎�<��uV�aa�noϟ��QR�����ܼ�%� }TZZϵ	$:�P� �9	 D�R���0���v����~���knS;��b��]|�������1a�d7��Cc|��R4Ԃ����G��򱧨e�y%0��d���bç�m
�-��������&z7K c�4b���3�H*8ӡ��r����Q7�+W�FTW� S���q�/n�|2����,��������q� �yFF�ی�q�y�z���.�Жu��#�����/��<��V̝��<�>��)�@��0Q%�0%�{��i��w���I��aj�g؇��̢�f���v�:�ƴ��;'�Ko-��.��/e�#'3���TC�
�\���Z>���1*��c��9�?�
�Nf/N|�2��Z�x��tR$v�'��EM�.-�9��Ң\7��CŁ��b�!A"@��KM�������?y2���j��]f!���DD����X4��a�J%W&��G@�1r!N�2;
LU�.z��v��OX��2�j�+��jddb�Ax�[ª�|}W7�TX��Q��Jx���E��x@�a��7�[l�M@�k���1	-x���Qҏ�^A��g� ���[��4u	>9U�?��oX�o�x����Q9��4u^6����	\����9��PK�,s��8��B3�]��Һ�e��Y�0ց�TnS�"�ؔ������q|-���'�/J���6]�&@��[$�sf�	JЌ@F��]��� L������akg�R*4�5���	�#�Y ^ �D��tg��)q�"P�����u�q/��u`�yp�g�����`�+���ˏ`Dި_�L�����P��慙Y�c���%P�#5Q���Dًh������h���Λs~�_GA2R����p]�OrC͞��tdk������ݦ�\Dkjj�����1�VϞ5V�<y�����L��-M�LbjjS���h����cq�� H. !T5���ڄ5@	���|=��M��� eحS/KI���e|?����t��WG>Ua�z$Q��Lͫ����&�Zf� ���F*�S�J�ms�oǈ�k3FB=����U��0 ĺ�~�Wq����>G���d(�����>%x~�>�	�L�&Y�
�� Y�#5��0tJ�/���._B"�����QR�5��}��vu6��i�g�-���'4�"��dXnecCr(Z���#��6?�U�	�b���`����^��i�S�$��NQ�M<�BS{b���t���?.����,�٫"��\�7�p��	rl�5�I��_�H� u���{��T > gi�l\_�܀<V�� �i@�h@�h~��P�Λ�� 6/f�%�%��6�w��VD_#c�
8�NM�,h�s	bN�t�-Q==7� j��;]J�ƢY$�����T���,���u]�a�� d޹��nm;U�=1!�G�����0H�gte��Md�,)9).-=���b�rH:U�ݺ��_��>{EaEA:�f��glf&��X��ơn���^�!a������y4IGŻ��+]�/>a���[=���/ŏ�b!���B�ZOL�Q|%���*��CHJ0_�J�h�w�UQ�2E�XBF��9�ZN:o���h���ޅ�߿��HV�k�OM�y���}42k&�F��ٔ귃2P�DB �Ld��˄�In�J4@�ҦU�^625���P��<(+������6� �b-�<|}���s_7��IZ����,?��c���^P����^��TvX۔�/�o�o��_���>~�B�`rn��N��h�6���� �#�w�U�Q����' h.�U�5*:Xri�� ãY=��N	Y^�(��#R� Y�Ȉq}�*� WXH��,�� l���&
�a "f��`��� ��z��`3���o߾Ex�֕M ��������_��q%�yO<y��Բ�] 2@��j�����a++��s�Y����m@y9ڊ�
tD����sZ�a9uH(H��Ľ��OzEi�y�h�b�c�Z!��u�j��}&�Ӡ�uD��Ec*1�'�E�Y�"fXo��r��R��ffe9;����_
��EsF��0c0���k�W�Z�@F]P SSS
�"p��j�7PPL,�Q��$�@>�yKH$�I�u����7�t7����￢���X�B�$���>{�_ݣ��C"����P��Y�#��J�Tu*B��i� %�1n��=Rj�'�@��5![c���|.���E�V�Qˋv��5_U��Q�\�ʚ[�5���;� �a�r��!�8"�1"��CE�DGWyz{�*p >.�����14k�I��~�%���#�;��������mݸ���&�@���1�VUu�&�]D{o�B������}vv�m�)f�^�\܍�zg4��a�e�|���b��������ݥ�*9��s�Aa��!*��z�
�J����`7o*x���yW�-� �K�hBh(�m�{es �#�{�~�P#��:K(r�3�E�
QE��B�U
�0<J;�������3�=W�{p��]�����Fr���K**H����ﴶ122
���G�A����Xb��5ו�ݮ��5wZj��[[��P�;HIE���� 8OVO*��à�����q.2E��ꌅ|p��>�jS�Y��3dv�\�3y$�%/�p���-P�~Q[)�z��ǘ�& 5��ԯw�n4���7��.��2��\�D�ݯik�{f~g�A���M�AC�$����Y>{��qٽ��f��v��-�v)G��{�������M�G8[[S��g�O�24,SZzG�u>���b��7EԜ^`!�:..�5Ů���-d�R�Qb�u�4b*+t����a���@:(Q��A�1��)b�/{?����¸N뚒�m-6�\������a�	��Ɔ��g|>~bwx]�]J����K�NDq�u�\Hb�x��\jG�� ��X_X~��X�߮c�J��`#*����n��h�WJ����d+Ɋ�N:0
�x�b "%�졻���T�7C~/�)ll4�Ѕ��s�ܙ)rd�z���"0X��|��Q4�~1
@�wAӨxZ.��< ��� ?�Wq����+$s!�@��{��l.���U䢸�$�����d�a�H�I4�l ���U_I}���%a/%�d �������xibn��t��g���=�Z������l��[�Aosr��n/�nA�p���u{�y�����-�э�h���\��5��B����/�y����4�{��&��V�9>�$-�8	p�� X�Y�{C�z�.5!@!OBd�/P0$���:�������'���b�}A�l4���4���v�`H�{��9�7[� ��T�� 1Y��rfX�D��8�9�o� ������1�R�(+;zo�7մ#��'�d����Ҡ�y7����ܺե9DHS�d���b.���&?+�$�sJ�;�g�
����jj�hCZZ*���ڀB��H\  ��\��?�=����z��z��b2 c��k�'�]E�C����dH��� �ygY3�0œ�v���hp �ᢈ���e���g�.��+�CENy����e�LJ۠�*�|��ue������!�)��Z3�і�>أ/���8)�˂7߾�W����8\X-+�,8�
�����X`��/6�T�SҎ�x⌌�#']Q�X�.ba���?���0�ǻ�&��3O����
��)U��SJ��ӝܮ<w��ڢޱԑGB�(Y�h<T�<$̪�]��oc='���䩔��~��6�",����H�{)O?��=�'��+�ͬ�Vl���u&@̓�-.^H��xp�?��B0�Z2[���ʛؕ������c�8R7�A�]�I2�J.��
'�G�T�YԎ%���'�hs�q���32"�
���;�5?Y��"��Ġ�T�d����{|; ���]�L=(��7�/���7�L�t��i�NO��7(;z�Cf�y��s Aк���L�t"f6TA�����2�E*����i7T<ծBa7�:���hq��龶��ћW��؆�nˌ8�wD��߄O�;ՇyeT(	Kx������k����_�8��Do��M��������Wb��?����;�vS�R6M�(,�C.�kp'��?�.�ך5���[+���֣#aqf�9�z�M*\!'77�,���S�-&�K�C����d���OH�6���>��b^����zǦFq����C��_��R�s��f�A2��+T�d����| ��dfib�����l��D@�dr�,���]�Z��W�9Z5����Gr?m�t���P�A��{e�Nkr���Zh����o�H<*���_�Aߘ�l�*���A  X����|�'��u����}D;�Ho��j��]��<�r[<�@MKK�M�/W�>/� �3���_��6]����g��D4(�����A�(�J=i�a���^�?e���,�a���~MS8σd��������Ө7��'("PS�ޡ'�q_A��p�,w�����<���]V 	!i����A����5��X�4ܠ��o��%�РC��ڪK�>o��	jb�;����M�ȺQ&W�&�����m�K�擗�����bT$��q++�?���^~A_�D�����}A��2�Vv��U6L�!�9g�Z�|9YX��yR��z��ˇ�::b�d�_.���iॿ��p�<�H���{�w��S@�:���.+�v;M,�~�\Nظ�0�s$��!��UN���&��u}�E�=�8HRM�U��B4�!w �uFrR2����o�G e_X��=!��6�V��Z��{�H)+��rzZ�իi��?�Ԉ����q%\�%�]$edځL� �[B�A����p�d��������r�{�Nf���e�.I��hL����G�I(��j���>���1�MBA�_̄����F�T]���bE1Ȥ�q��>gı�ˈ�7\+ڨO���@��[R�_�z�r<�w�sUmN���Ag��|^�:- ���d��B7�>O�?UI��X9��;�Ź�t������
:1y�[Vf�=�/��q�n�r,ad�+�����Z�������$�m���D{���Y�˷�_C[�|6.|� �d��޼�K�	�&n[cK����3.(�
h?`9�t.P��*Ε<�,��x�`ÿ|��,�^y��P5�GN���s�Ms�����A�7ڡ�OZի�p/e���)�a2c>��3V���j\�:q!H�:E�埰V8-�� � ��z���'��d��E]uu�}��Z�~��h:t�Y��Xbjj�Q��e�33w٩}�y��b[�˿��<}z�P�,+ͩ�]%�C�k�76����zl�V��:��� �����ꇦ��Ŧ߶�=8����j�A��Ukv��
ex�)�<���]��n,U���
i�@V�Fӆ�sv%c�{���,E�|H�x6��)�l����( ��!�#�ҟ���D��n��>�<a�v���7�Q����w���2�;h#=�[�?�-��h�*�K�������T�7���\�Z}}}�L���6����1�6�KGǫy�%G^�/ww�A�C��[�gϨ�,K���쏏�x��!Si�[�q���E��oH3����X
Fh��j�A�k��є��~{Mc,�<�<AE�|ԟT���/7�l�'��i�d6���n�]�Do5M��L���?�ȉQ�y���wx�|d�}�Hd�\�]�� �ey����*��y^Z��4��b��]�%�e��Q)����aL���{�SY?�5�B2+9���w���}�إ2u��Ʊ��V�=�����z��Ւ_��6m��.m�sq������l@楥� U�Y*�WW�/. ��W)�5p�鱥�mBV�۝���d�F����.3T�׽�IE�(������7��|��D"GE�.����xɫ�Wc�ZO�Y��%@;H��̀����R;Q������Ap�
�&&7@u>8��`e�G���쨏4��pZx��Z��e������P R-�ˏa=��RL��kC�`�Gp��b��R|������̏3��-+�(f��VV�=��11�V;�
mڥ�NA7�B���8(1`�@�-7���jRl~�F�&_�R����R`'�O��vE��	�AL�E5����� � �F\��(M��q��7A���f�`��DL?a���]���r���Ce��ޅ����؞��饋��,��g�8�_ �_�я:-�����[�>�4�ǀ�%<{aw����e���Mc�2 � �t�����_�ܹ���zw?�;�;���T�k�QiDx��+޿ק����ո�|��L쐀W���-��b�����gg2�_��
��u!U�z�7���hv�~��q�O����+�~V=Qs*+.�:R�R��t�������CP�+�/埇�;��g]c�+�l3�-��6�w,�Ot�.�$P�77J�Mp��YT`Ra���!SԾn�졁��0�t�\��g��\�Lߵ�*���g�hb�l���x��j�!������ޞoU0?7�2NS]y-َ�oc:����d��������gR,��9�-lm����_�n��w�1p���	1��Y47Z��sjj��P3�֨���VKojf���_��1��[ʠ�a#���,�J�!�Z�X�꣊!���"��Gʈ��S��e�7����*���KM�����b�kh�����i�/3%eJ���>��ۀ���{Ǖ�шh7��� ��M��8�L�Ԕu��<'j���}���L�G��D���ٶ����/��?��O>��W^]_�=U�R�]պ �v&.����W��������bm��=� H	�i)�s�0"���~�=��^�2vqu�HU�ՁFuZ���{�i>��_^�p�a������-�5�T%*��5_$�|��[��px��[gj��k�`���!*3޼�H����2��тJPE �3޾�9J�r��˂��0/(�<%�ϛC�
p~���^6���:�\�L�eM9l�n��H����>A{+7����QT��F��l\�����h�h kfN�*���^��?''E����y"
����Lk�V��~	9-�4:�3�B$�h� ��Iz3C�;q`���
@��}�l���C��b`)�'Εչ^=���2y�.��v@�7�B���*%���D"�k����EN��n���^h <y�U�X�Q�ܢ�Dux�44T�N�6�,�Kf�eB�pA ���yՆ?9���p�0F�"�pf�;�
:w��\����UX�,Z��2��x�d���|] ���?;y��{?@hC�)⿺$�%���C��ޮ��O
Q9ߓ��͔���Q~��dw�-!)a���:h )촮�X�	=>�� B�Y_��]78c�O����Ԥ�Lv�"~��͸ny�#�\�ɔ_�is��oQ��^R�%�+���/����GT��/� �ɇ��P%g}!7��A�`�V�K��N�P*^��O�i)/CL�-$�FM�ݹ5<8�Ü���n@U,AJVS[{��-��J���
�D�9�}�v�vǁ0�Q�H��5)��\_'� p�\J0��=Ϭ)q(��
�{�@�$@ہ�8)���d�	�����9P8%e�F�59��w�G!�����������v�|ȇ9C���� w�FS!R��1
������tt�*�����옟o~��Xˇ�Hˊ�n3)���)v���d���vw4	wv�Ǭe�K���z�162̿���ՙw�q�P(h���̮.�������@v��k��cuc)�^���<9�~L�o �(�P�'����؋R��X0[��5A���\�����2Kо�L٨����6O�5W�%r��Q��w�A�e<�rswV��ꋲ|����b` ���y�t��i��G2��R2����\��E��<�:���1�>�L�j�x>�x���s��sCFN� �}�q��G@6�5�����	{�u熄�S�v����VW�X�m�{2 �`mk�T2k�f�F�+��"B}ȁx{��UÃ�Cd��� dq�Z��/q��:�q�A�S���t�޸B Τ��s"�29�:!-d�
,}�u�7Ksuo��̙f�����0��S#/������'��H���
���xi��	d�z��X[�0t���<���12�����1D����M(��6p �Qm
������&S��e��a�yXN`����s��&AJ����L���Vf��W#�cВ���|i)hkt������Nn˟�o�G~N/d���9=O���Z��^�\ĘY�W��t�r ^��W�A��/:9�:���\P�}�D���m@�Y$o ␉��7s�c��� d	j�&U�O������,�Y�C>�]� �?��RSS��=qIX�犘��5᳏��g�C����ie,0/S��-�w�0�F�EC���О�o��o�UO�&�;)t�6���.�΢,.�sm�73�O�ې��'#��M��1��sUv�gb���@��;�����zpy7���ȫ��6h�1;!zPR鴂�΄dBH�����&���	-��K�V��_J[�Q�d�E�o���(��-�5A-�->�5!kO{�Z���/4���/t��d�ok�,h?��������Vܿ�p��J�^�zk�E��[[��������>D.
�fFF��!/��*Y��ch�Z���GI@���|3a��ܜS�il����>��g������&���hY��>)������34N;�U)�:�V��v[>�ܾ�HK߀�iS�7�-{X�iH����\�@�8K��ѡ��7)��Ҁ	�}7AN]���b������V�F�K���Ž{�z:-�����X[_�1���kfF�PwEK��/��U�8[��OQP >ǚEq��H�ԅ�9��I���X
}���D��d>" �1J�m�0��@���;������uR2�6���Ҕ}[�йq�g��29td�@�����9D��nSn���1�<�Y;%�(�n�	�b��;�q����̜N�g�eN���!`X�R����ѳ2����ii/��V��5�C��y�՛_)���H|�v�ʠ(��f�*�ץ]�E��w�h�0	�<$2U,h[��Y�=���,+�=zKԕ|�V|�妩��=��ɵ=��n��+*�*4�9�̄��o�Ǎ�ߑ�&���i�+��v�}�]��Ɔ睕���nϥ~�OO�����3̄�Q�\}w<����$Tv������QfF���{d&3�C:!������qp̬����~�����qz���z]�s��uߗA*Î_S�2�͝V)��s :G���	Co; ��x���ڸ�� �ǫ�w��y�H'�N�-E�с�#�-�*K�z�=�sʞ���s��N����"X��MOs��U��%YA�
����-��?�9�@׏b섳�:��!��Y�h��{��.V)U���>��T��˭����B�J�	�^���E�_�V�e|�W��=�����G; ��'-䵯�r����.!�3k�r��������Y�vt̼��R��y������/��,vq�{�sT�_CDY�a���è���HVF�����DD� e&`(Pd4$���n``�^W�����Xoq)�*���,+G��wO�D 
Ϝ�FZ+20 ��|h�CS{�G��%��?��|��P�H`��v07�����e�`��y�q�z���<* x|-j'����<��aWWW`�0�78s\*G]%�\�3]%ze~�T�ԉ�f��5��WG�W�z4�.�w7cZA�����c<�Mp��b���9��U(��N�b���������,���/2����?���"�l,�O �L��C ��(��T5&�z��$01����$��Lֹ�(��z:���>�����O��+&;^���'t�d�hbPӗ�6G
�d����H�E���N~�%�<���K����ڳF�s������݅_�A� �E�3�c٢�ed�����[ncS .�ۡH�`�F��D�yD��,X���@�����Ig��=�@�d��߆,�ѯ
4l��6�0v�G��:�ׯ%�uӳ�Z��ǿ�ml�����=��4+���4Ӡ_�r.�{ֹ.�r,��Q�Mi���D���8�VO`�������d)��JM�;��ݯ�W����h|��<3��o�Wֽ���a� �1E�ܼN9\N��0=6�(�����WE/4��]/�]	���f��Oc����p*�.Kʚ�Z��;J)f�>5�jl5|��s��p�mb�sJ@�s��yO(��/�qwR~"O��ʵ��t���I0[�����N�M��B�EDkɩp����j��;lji�
j��z��eceDZ�ԭ�Z6�$�t�{�\�Mu�Wl�^�{x���p#�cq��JI'�������A�2�<Ԣ�$��nݐ>ZIʘ���]n���k�*���ª+��S��CC�f���M���߽k������������#�1`��w�F|-9d)��k�kR��~ڻ�]Ž,w����F�S��C��q������Q�S5��� �k�'�e��hnȾ�a�"��E���'�o�k�����=�sR�a�Z�ǥ���b�g  ���mY��͡� ]��s����p=�O��+��C##�h�FJ4�N�s�K��'���:�4�u�me�DV�7�Ȕ�0�C����@	�������֒�Q5O!ͭ�?,K�n�9e:(�jE)��D�nLq�g�J���q�m��|�|�/����S���/�#a��;W1<:j9;�hE5}>s�>u��oJ��Hx�M�%	��Y
�]_�VY��ATy��8d�]���ZT���sV*���c����\��(�y��y�!x5�;��<�_�+&0HeW��y\vF[
�'^�&Y���ϫgߌ�O�'�Ϗ�U������Ĵ��F
]�W3�Ǥut�b��)_�'@�U��:�4퀽����Z�D�$9t�HʣK@����5�rNE����-7��.jj�VnF?W��2^�����Y��2�v���c�r��e���~:�\�6.��NA���|��٘;��c\�Z�z��AHh��7r���tj�Y�s�.��:�/��#�n���Z�� ���V����=&2_)P��뷉�!��C¤ �b������}'�Jy~�����*?�VTN:n�>���C��8~�%C�)����(oK,�������G
;�F�����%%J�����D���R z���R������-5E@�;H�+FHD���GG�a*-}6����a�`����P3Ƕ����UT�Dw��_�φ�$��x�p��,��x�Ĕ���vg��;/>��`۠��>��Q��\ZUh���w=;�غP��Cj)����w�����i�_��/��!��b�̒\u*�w,ohh��G��am�<3Z��̌u�<>���W(�jf���%*�!z���������+�^�O�&e����O����h���}R�k��QB���+ޒ+ޝ�������GHG�e��c�m/Q�� �^��ݽ(��%�g�ߙ��K��F��t��i����J�Zb��ƀ�^����j 9s�DJ'S���[�Ul�����;Z�ij@��rБ��7�
��������yyfQ�� d.)����s�����ܰ��u('�����9�r� ��D�=M��wW�ր�C���N���@P����`�������e	��C@&-���F���"���^TD�e�)�_g�'�F�9�ח�|����؃W��i�P������#���]^''d�̢�Z�^����]ԟ�an�OPR�� Ds�������ŏ�O
�O}�1P��j��E�;8\[���^{��iG$\C��/5a<�-˻�J��\ިQE1�{�1�����FC�� �fB��?�Rm��~��U��_�wׂ4<�,-8�Qt2KP[�ݻ���Ǜ�y-��j֮�7D��B�Ot��į��D#jk�Uy���E$'�=T����\�zqZ\����j/+Z?A��<k�n�p�9kr��8��ߝ@�Jw���R�ՌM{JL{�M��O���v����J'����is�\��������ݪ�rrbl)T�����;��=�<�ۨ�q�).k| ~����(!��E��=�����Ef�뛘���/7h��}A"��եb���j��'X�(D�:~-2��o��[v����"q�ؙ)�r��I.#��{}}���O��3^���B�~ �KV�&���V�y�0�upw�F � ��+�N�����]^����7#�`JE5�� ��W�KV��\l"^�Aj���r�ו2���b���z�� `�̤M/r���pE�4�j�U/����>a]���6[f:;��ͤ����KM��o���hxX��������2����9Y�;:����T���=;t{��S�����:��9�ǥ������G��\�] ���I~֭hJ�H)s؃ؙn�ݨD�}P�{�)c��ta������l�ݳ���;��{�AK��Nv�41͘��ഇ�<�>�C̈́�%��Tڝ��]<Ƿ9�6���SL�Mm��e<�z������f%�h���A�^�^pչ�~��$�����aj%�V� h�8�v^����խ����Р����|�.�8��d='~ [)�a
d&�7ʇ�f67M:%� ��XT�}q<m�?�	r���j�w��Ϗp����Oaj*��e��D�}�e����?����|q�~�	oڕҥ�5�_��; ҳ������,#��A{Hsf'����\#� p�L�߇�S�}^��]���{�S�9�,L����#�HX<)?$;�QJl�K���fJ�(�|��x@�,�.��_���뿥&����o�8I[�$�2�5�,��E"���48���t�����!�k�������N�X5�^=�K�b֑���V�G��_��g��yeO��Hr�:ryO�m��6���Y��j��;��|����g���+W���Fi��v�&�����E풒N�!���\k��gb��&�7�ꂃ/dkڎr�OO7.��$��╦rrp�5G %��O�*Zo�d���=�A�s�@�F{Z�}�T���㈏RR��Ώ��jν;_�R	#��t�����%�/����)�d~��fNN��n����>16��M�<; %f..DYd���=�E�����&�#��K��H+'���{C� Z|4�AA5.�S��O��+y�P���Ž{�)\�f�A�d����U���	4n��BJ��Lx���EeX�7�~PAԊ!�5�}���	(+P!�J���R��f/�fD<)$q���]5,����6'k�����л������G7ڞ���x�]	��XB/��3xI�?��V�O}�=��I�W-¶��ϟ-K�q�aI�e؟W,uu�c��g��ޑè�:�oN�Ţ��d?W�po��''u����ޙ��B���!�s���%h��4NL��%Le�w��� �X
|DP�R�6���+�K����g�o��V���$������s���8��m0)+9C���
3|�:@OX��Q�J�	�y9���ޅ�I�l_J�NB�kb�FAƦ���v�܀��~q���,Fߧg6	��b#F�u�B��BW���wg*{�#��H�(��x�9�!q�dnD��|h�݀��e�mtTDuÉ姽��.�������$���tJ���`����uꚩ�Օ�EZ� �O/��4Nt~3y:��K�e�0�	��̐3,���Y]'������S��L��D���Ү���'�
���YY���i��N�ȿ|�Ni�_�",)�8O�]\Kt[���G �:~��{�<�B�9�(�*W����@��Z�)}����Y�|�gKo H%'��Po�Vґ�J�$j�{Jdm�(è�L�˦�T�><a�9닅U��Q�EF����޽[�����m_Mc���S;�qеpܿ{��w�� F7��Q^�Zw�j�I�ϟ��&s��P�k}O{����`�rT�=y��J��'��`�X"PDiC��FEE�}^��[(ޜ�M�	�$�ɺ\��>��A�Fh3�\�����u�ե��.*����3�/UL�[F���T/�� �U씁Wj�bWW�So�.|�7�Y��x�E\Q���1DǞ�U����ɑ���D�Y�$yt�q��r�)t.Te�Rﳿ>�6)�	�y��2��\����V�.zջ�!¹��_C����G��N�u�zc<�ؚ�:B*#~1�D���u�4��ܛ޸���,y&t�v����H ��Ԋ��Fj��UK��M8/��m��z��P�r�f⇶ ���ڳ	���>V����^�z���Pm�U3[��0�����f�7�û�1�(�jNr��G\�fC�͎ �z	C�?�����dZ~������=3#o�am���vu���� A��ϟ��ǜ���l�9�3���751Qc���h�}Ë������.	f��^�WK�X*�r�Slp2Ĳ��4�җv�k��4.|�U�w0���R�	m�s��E����2M�7�<�^��e�xZ��YW��O���������	�	�Z��:7/��M��R@:���ȫ���0/��s�*� ����\�(W�= ��k3��t-�wW�FD�% v6����M#�\;~)�/MHٜ˂[7�Br ��I�G��bݩ���Γ���X44s�wה�|w�q0]��]h����\Z����:`�7�g��Q�y�<a��:�WVW7;`����5�Y]ݸw��1�?�<�\c�T�i��K[������P�RE嵐�}|�V���F�J�`*đ����XRSSe����B��q�=Gy���߻׌J���"$�^�%c��gT�k�Ɯޢ��S�YY9�db�eS��JTy]W/��
�����ꪗ3ˇ��~GQM>�+�g&������!��	�1�/Qy�B���h��'47�xRl)�NMo��5��U#�m,�� O[׏��_��M*�P�S� ���b�f��'������hs�3�Z"_�[H�H�M{z��JD��e��D����K�0����fA1!Q��4?/J�(X"y��"W�כ����8����w��t��s�WK�Ͷ��p���^ꋫv!t�� J����H̀|���g�3��&O��ʪ^�}e��8謋�(��J��w��2������ �m�[��k4������$�~�@m�Eb��:;�^~�M_��m��]���畒j1 �E/�a"���5�����c{�tLB��#9S�A�����MDX��JKd�θm;H��Ꚍ� ��o���BL��\��ۯ���ѵ
=��х��!'�UJ�n�M��%f��#pK�b	3�źF���$�4��EF����j����L7#��_�+��Y��Y��2C�^�23�zU 	��HB�t*jx|\N��������ȋh�Hmz��lQ���d� 01[e�SS[�u�O�ҩh�S��[X��ݞ�6�7Vw�9XA@�5y��������1@&�����,��S�+���1d��S_��W�#1�\�0�� _��#E:Br���Ն���W�Q[�h�P�\sy�C}������d$��2Ԥ�z%z����5%7���
 ^tRUR�����Գ���J�g�J��G��1��
���ۻ[�O�;N��������MM���KM}������V;~�Ș#�nm�2����	��qBE4��c��=��3��bFڅ����,�g��v�2Y[[�"+��W�.w��_r�S��J	3��Y�H�?0V[9QkD�>�l�ܤ�_�����kp8CF-.��YW�����ux����"�T�Wr e�W*�}z4���3�=-�z���0���-�gj�&�aT*:���*^`�;�g��E~�E�1�J�:�$���s������"��A���p��KW�r�ХP�?�,_n0ps��'�F�-�1u�G{N�-U�d��}Y��2����"�춸.4�����,d�+
/��/2�H���-z#�����������4s����4��d�/.u< ՚�9�-ѫd�>��j%�Wv��Jr?]�8D��2��+
׺g7͂N����d�m`j���܄
������@�����á�1�d�`ɉ����Kk|����ϝ�ɀ� @9����9
����f����j��2���_�T��ԍoFΨ�^�<41��%[�M����e��8E�t~�p�H�Đ'1�2c����(���	^����ش
�(��Y'm����@�,�W����$�/6���:��KY�e{!��#f6N�sX���ު��us�4������/l��T���@w�1R�;Ȏ��CI����k�8*+zc�I���Ӵ�U�/��(�a�L�K��b�nii�x�L���q�I��f����_�:�j���W�}M��,�K�u���� 7<�~Kk����Y޽{WS�4K=��S�bvM�?���eS"��π[�	�Nr;��#z]�}y�k�u{����k�Y�,���VF|Q�&5wف*P*���0�Y�#�QGu(�(p,p��ͥ:�$��Q�u�C������sl)@w�T��S���U�1A\W:K+svυ����iW3TŽ? \�q�����g��L��ל;��j��E@�[f�Е�]s��
�@ƕW�W��E��{{{�Tz��ַ�����Ls( #Y>�P�\��Y.f��;xH\ZZI!_92�,�����j����Ο1%So���8̒� ]�I9h:K% �djo  y�*���qH�����̄�?�W��L�������S�M���E��x�����a�[<Xu������,����/�lF�䙡���F�pz��*޷�ٷdԸ�HL���k���� ����#}�)R����|���tu�wP��ѕ���⧾g�8�v
z�Ƞ�%H�ߤ4��Z880���{ׇ��[nVY�o ���J��8^�2�444�^�VX��޺k@ I��6U�� �_{���0)�n��
3x�R�,N�)�}F�Hr�TI���Dھ�W(]�b�XϚ�p��S�Ì|v�נ�Y��� #0�zH�T�H�P�eXɁ^P� 4
{�OPr��T��a�zc@�Vx��P�k���Y#��seďZp��w��#1ji{�S�=�AޓrAz���]�ior������`*�$��w��|Ũ�s*ڸ�~ꏗ��f`U�P���j2����g��kD��@*�8�Rș����H�Iw:YY]y�W�d隴EeAL����AH���.�{4���Y�o��RӞ���>Ɇ��5�{��$�X+e�ue�<Jo��w�w�UDop	����_��n�L��VN�p0�0x�`"/
o�7,ႩD��6�Z��$Mm�&*���:�����7�� G��n��t����l��pBҊ!�������0N�bڪ�1J�BI�o�l�R��{�gǾ��I?>��_��l�w��]]���f]]`G�N�n�}#�Z�8E�23�<�Ia9<�Eˇ�i��U���U"��ݎ�\Z�l� ���QB���z�������X ��
��`ޓ����S<Q11v�����99L!-�R���cb����z�^1���E�s��������=�U�l�\��ϟ�����(���t���r�y��3��~(�phg͜��A�O:�Q
9��]T%��
O���mr�Q�E}��E�m��":�4��B0U�:#@��_�Y�yOB�/��i�^
��� ���u��
�#n{�������/�P$�%QWW���,x������YρϚ��ο�#:[#�W~zpB�2{�C������go/|�6&��m�w/�X�Ei����b{4_�S׹�qlL����-5����cY \0�O_ }��zqQ�TT�w*.v ���.7�vhN������89�K%B��qr%��m?�����0C��8Ӹ�X���F��g=���������) �[���	�$2�j�&(���%!
�b��}	ޏ���~? S���0����B���'c��Ն���\�9��l�Ed�M��B��4��Q��V��9��B��.�Doy~�
8=�M��\ڳ��a��$D��x�W}�������45>'�#�kU���j�I��V J�"oQ7���𦚓ఔ���Q	&��dM�w��Ltʟ��4M�̌<����Lq$^6t�ތ66��3�c���j�
��u���¢w�&�բ��]�v��,@������Xh��-�]��O�c�K�(��&OB�ë ���@�E�j��R��כ�ƺyO��h"sx҆����^�\={Y�T-��5�T�$	�_��wY;�t��o>L�-�9�+O����.gȁ��v�=/*'�<��겊?:�z�uP�&��v�6�4mv�vb�t Pϖ���i�����ʥu͂��1��|�_��I�6ϊu�kjP�L1�����m--3}��	hJ��3�%�s �w�û��kLSAp=	aׂ(�&~��S@��=�����j&�2�.�4��P`00((E�U�Ȳ@KFv l~,�]��,u�n�IP���/̵�f�z6�� �:K+A��)���,���S�C}):g���;�{ar�ߌ�����wU�q���⠒ccjܡ�sB��
�cw2����a����m�d�g����wt�b���1O������y�=~�X���.�E�z:��0A�iW�t���X�UGA��Oxq�u����s�����5��#�@$991���.��R��&Vђ� ɡh�w�#�J	������X����(c����@#j�q���[�:�k5ת�W[k *�."���i���(�2Lb`��1v9�Q{D��=�J��W7}��h[����4���)Æ��Y�$%{@W	���/ kUV�����\;�8�sz�$H�S�M���)a�� n9ӳ�?c��,���a��4�ǭ�/ƤN}��)Y޺����'�f7X��r�ۣ��mIIg���]?�^����ҿ���dT�IY�M���Ʌ��n�C�ǲ����z�&\���C'�������	�"�Ȥl�ϟ�qq�!���甾/@�R�Q�mQ�eW��b��nTc뼆[��_��y�o�`�{-ӫ�s^/��)�X�A�æ��������r�έ˓�c��o�Js���HZV��]����P�X"��� �\q�U:A�3亂��8�����u`I�c�%�T��þU/ɚ]�F���1��ͻ�2��M�{�o�OFWi�N�M���c���rp0�8�@}g��� Â��UJ��R��^�����G�<J��Jɡ�K�rN��Vt�������]��[��JF;-��B�f�KK��UI'������^�Lgw������#:�-�A���4���p���E��#�=y�qs#�V�jƦw��{�p��Q �]��t󼜸uje���|qz���%i��NM�oh9]^+X�M�91��H�J�d4�n����Fδ�J��
5�j�d��K�?�	Ϸ�I{�w����8ch4��!N�F�f���m%#�&�h���%�.t0�.�_^fL�%G��/G{gBA�	�ĉ��G#PE�V���e�/55����F.іBỻ���$�|./i	�ј�;���˳EٵU`RD͓vR�q����	ҹ��('�"���;�	%P�|�g鉰��V��+���+���.� �+5Ռ3��7�{2������?}�/q&��]s�R�!��o�*è�@��@7���p����]�`.}�!�|m�M����7#D����B�C�4W�+ot��,VT	҃��K�����vκ}.qN��KJx1`7�,k�;�ag]1W�5@:~o���o�˝!�#�ց���@'m�:������%P���]c	�+Pk�T����MMh�j�d��;wLE蓭�+,R�/{��\�{i��{�6�{�%�"V782X@Ƶ?����Y��p�H�pNp�5�*���Һ�;�P�*V�9�=���'��z�+���\�{P���FQ��4�W���J��f�8�\���*[�jÍ���RiC�Ld�Y��1��ɔ�'A�h[�q��hԜ\v�؉�J���d|���vSQ����0x����l/I�J�'�� �7���BC˚1�X�=�Ajym-���F|��E�	(k�A�����F��zpdr���R�L�?������S0�q��(��͂t�R� 	�w��v��6*�ͬߦ��c'��RȎ:��˱;mh��
�*�DF��C�̓�^����"[5�+Lp۵t�=�����beu{�j����o�r)��@\�D����T��[�,��>	(~�{�2?2�$hR왨/]H�Iy��O�����V@
cؙ��������yD�G�,N��
�A�u��)@H�n�R�M�35���kE9_RI�R^n�b{kuL�'�h^+tu�+C�0貚�565̗���-R<@߃N~D���6v��Y��A}����u�N��hZ�L�3̋�( A�54�|��;���x����r~�QVY�]5���h-[��IǴ+�� ����'Ag�0Nbt$	(+h�f������-��:���?�	1?H���:��I�Fs%�։�޽�9���y�5�B�<�0���o�l�ۜY�c�1�_������C`�;	v_�d��	�b���:L����N<~fd���h^+��K>~~���1������d��}GU������<�
�0T�А�,���ɑO���a9����5�<�-��39F
i�?�Mf��C\J�D��'���/��7h�/���"NuǄ)��M�gĔ����}��	���MӮM��;��d��II"��K�P�4���'#~"�TJ��Cz�`���]�ڎt�q�tU�,b�>/�jÞ|O��&eD� A���J��c�J��9����1Hd�f�D�vG9�9��@B�F����ꢥ�g�m�/e�bT�ΌD4��|(;?/"}�7'�K�*�>'�O�
��ݭ
ޮY���U�5�]]_�G��u��
���:�hRV.�ǡ����O�I'�IF%�� KJV�*����I��=aq�� �JCC����
�>�vzۿ{�b�$.���ϯ��/x�@n�!z9��"'ϼ��:�|���)����բ_���)�a�aT���:gAm+ek��/��>j-��}�͆L�����Z�EP4h�I*�<3�t�2�7�)�K��?|����)���,4,5r�I�lÒ��.��J'�d��k�/d����A>�ABJ&�(��u���oJ4t>��r�S��-�ۺp`�

��l��Et�\�mcly��OO�+��--��?k`xηI/2>A�*s!�?W����,pd�w ��%��ea;����`��@�_	�����R�z��v0�'�2�g��7 �9@�����}��\t�aI����=4�w�L�Z�)tۭU=%lk$�:giR�r�t����Q��^���� ��~M�?N�J@TM�=P����N���)9�`�2�J�/�E��|_��*�HU��*ް�H����ߜu�=��W���}��K�AH�D�ɓ��O��{��"n�Ѕ6N/f�G��ԍ�\�_AۯC̬2@(��S+
������!㳲
 g�~��ʀ�;A����M���w<�֠y� ����$ؽ͙vJh�ʯ����zƑ���mYIO}��E߆��ҟ>⺊f6�=�B=w��O���Ks�7K�PՆ�'����\�j���lEt�Q\����eۚg���L��K���i-t�u89��o^'gKC���'��QhR��L]>�VI��Q#��s��*����Y���p���]ÊlYod���q2�oQ�=e8�ol�i�������]"kxt�fI7��nm��lF������D�ڴ�F���mKSi�}���rZ�,+�{�� 6���]jm]]���Z�{�Ғ�н���������E1���=����������̓���&����>�8nLQV5��4⿊�ȿ����ڻ��	_������'0��fQF�(l�e�=4`j;�|�2 _�L��\u��V��7�`��?ۙ_5,#���GK��i`>����nK�!S}�
���~��3f�Uuu
�-jjjb�g@Kr�L���N���?t�o��F$��A۞��u̹�����&��X�3�QMe�75=���3ڜ�E����=7�Y4��=<���Ws�򂐑��{��)"{����^:�ׁ���.�K"r��1��O�
�\�U���\F�S�eXU���Ǵ�����sRV����X�ձO�ֈ����I7ޔ+I����D�^��5ⷱ:l4,���q�b˯��-������ӛ��v��f=%ж�}˻�%�r�6�.�2_&�-�JZ4������Y(�%v�4� �5�)ʰs����* ���v d��!���H���_�u򵡎����芵��5�k@@��uk�I����@�O�����a����B/@�0��f�q.r?v���y�L��Ռw��L0��?{�����5DTV�r�'Zb`g����&�uW���Y҆��/����Ra�Ѷ��9tx�� Y�p0��hlP�}0,}�&���}:D��+`�̼H� p��l41𡃀  (�O��8�u�(Zߨ(*J*]>���u�؝k;��Z����jP'���u7��殪ި��>���Q�1���QA�9�ތd�Oہ��[�y�i8�%��g�ԯ�*�˟��*�b�~õ�~v���O��#a���%�~7��^Myt�)���	��h��Z��
�h��rt@�&��<iUO�����K���f�\A��us6���e�r�)����0hG�R��EY�}���
��)�[=n�9�Pr��ۮL=�-�QKS�P/U����������}|Y2�z�4��5�\����jG���S.��э� o�:��ù;}�ޝ �:<$�R���3fWɭ���~�tlmQ�m����{M�]{{$	|�w%���7< �~|��"����薋n��1�7����� EL�h��}utn.�@@:��O���G]]s	V���O�� ;��=w�6��XwO�X��@���3U�=�o0?&��A�r��x@�v[�o�p3�f��bgE&U��$(�TE�"@�E�Ղ�Ńm?~�Sc�x �5_-��HlN"�Ư���tLQB�R��)J2�gv��L���y~����nD��Z�����;q���Div�9Jd)I:ksf+p����131���	Sɳ��Ŭ�9����6��R�����)O2��B#~���{�݊G�k��Y�6��!M-�=�,��/*��n�7�Q��J�t6z⵭p���c�=��ҏι8Gռ�i8T?��J	�ȰVφTpM�>��!�
�<[L�!��>)|�t>�
	��fR�پU�ioU��@��ظ�:Z�b�@�ʦ�����B�,L�K@�RC��H_� F�F`߼�腓�oK�2f�yB�Ԏj��/�w�SJɿ ����9<WD�j��"�镕�|�7fa��^(k�V�/��$%z�|K�	 �DEEo���tY
:��%#�Y߳��"%g�k�s@��=��OO_��K��Hr�"p̀���L�]6)s�d7*���D.��n��&����DD�eZ@G��3V�mK��<˖���~�Y_��C<��P�˺2sXF�i`n_�n/�E��5�~���̤���zh�D�b��������#�2ktڭK�9�Op�+4��^�
���r�B���u����o�ju���a�Bi`e����C�����,�U�=pl��]��b����8�<:��.(%��kk���3ZP��d�Ak��
�Ά����X5KY�������S���;9�C���%^�+6�F��P[�̓�X��� ���j:�׻-�$* ���'�(��e��� r�����B���Լi����Tl��Z(�viD�Mz�\���,ʉP����vtX.�'����Ϡ�����4�r��н� ��w��xJ�E�?;_��č-@{�{���=]Yo�!"�Y�yw���}�o,���1��1��� m3Y�ux��}֡F��u��7q&�����1�FcU���y�kk_�ݾM�u�1q�87����«Ԋ�L,��O���x�2�E�O��PA��EYA��6�6!�r��2��|7��K8iѕdN ε~b�/0uW��ڦ/~ʣ�n����a�I��\�����8�L��f�^��Ȳ���tx��6���1����,��6$ض���D͝.fԀ'!W�/0�xS���bY�[<
$8�a�����سT����fM1�E�2l�������
;K0���B\#���B�`��끈|����
G�{��+B�����O.;��X޼�-sTV�u]�eyt��κRh�ӕ�') �P���r�"T����DD�]�}^�*��l3.�k��Aj�fxH���5�2��J�>�d��=�G�!r�g=̗��E^��~�	�Έ0O�0�ZU��]�M����؊¿���k��\��I.��8Ĥ,�W��pa��EOB!�&�������0kP5~Q�iJ���w� �7�C�����G� ?s���Ɵno��;&L��ǎPo�w 6ؠ���(��G�
;�˩DKh����3~5�zxx�zU��N�M�]~�%���~�*W[�m�JRx܎���F�u��)�k�h��@~�u�qp<f��z�[S�8:y��
 �D/����AZ�/ȺD�
�T+��0�T����9+�V���fP�N���!(�+N�޿��wA�+�b��%Y�Zot4������uN
bC�k9Д��v��[N�q������mTuAٔ�s�����tz#<F	����V�<ޡ�!5F�0���ɹ�vA��o�E/�̂�ɳȸGԢ���˳B�� ��~h)��#%�b������F2"Y�
�1�_��_��w����Sʱ�{�����U	C/�>��^Z��F��e�B�{n=��0h��=<9��ZŃ}KU��|Hr_���P�S�Ǳ� <4w���(��i�>�.��V���1H�4Tx�t`��VX@R�je�;H�t�F��J@���ɓ�Jd}�./�P�3�eRȃD�>ϧfݓ;^�g�8I/s�e#U|	���j��}cbbRi�a�<���)jA�#�OO��^k6��al��璒�}K��SU�V�b���g���7VF�Rari[�R�Ƿ7���lI�>�Ft��J�C��/&�G��׾�<d�;���vb��;����E#�9h[@��Xb�A��3�./I���� T#�����.��'M�@ٚ����#�Ts��ۦ���s�`�K���y>�$P���F�Ӛ�7\�:ʜ�@疞6iH�_�W{�)�L�e��^��j���X憢�s�"�V�X<d[���GlTSӞR���w�� .�%���e@�_k�J��\]���M��J�,��ʱo3�,���H)�?�[|�P��&&!����s5y@f�$�#��U��T�S�X�$�3�䣨���?�}  �EL�N��\�����������9�KA�ޭʲ��
�A��|K�<�v&�t�u rY�j�� Do]Y����ir��(|�_u�I}?�ѭ�CF>pN�]avě���	'.���7���/uJr���TY�L�xf	�db����z�2l�����O:���L�4*5P�Pkg��6oEE]�����X�2+B3+�Q?؜L쬷����S�$44��p �O��	^�@#���ϼs8 Z����&�ս�||J�S[{�[m=�$W�]���5�㣩����@���H���1nZ��H��HyP:��E����jH�	��1'a�c2�K������ t�k�P�\U��U��6�:��#����z�^v�3#fSD2P��7�.�P�?��� ��S;�?C�C��KM}̓B�5:��I�/�|h�jWϝq ��S���@I�{qs�߻��j�����cwL���/��܊Z�����ɧ|4@�^m���>�v�!{���m9���w��w�USJH X�|�A Kޓ��56Q=�H�$��ԙ �0�.�<���]��@L�m䵋�� ��U�3��@mZ�UA���{���eM:��w��XK�Nb_-A�F�X[ձ�����aB�G\�#MC�_�іע����t��<b��|*�;!|�|	��!�\����|��؀VI�)"=<�JCN���P>36�������VB0T��ms�fy�ƹ���9{�Za��8S��V�\�W�zh�Oc���ny�	�ɺkqx�	9���
�sv�H[袡���c�	g�2Sd��&e;%zx��ز�^��t?@��S揫8�k��
h{�ڔ� �$t�0��S�1���.��w �@�
�RO�
�c��4BfP Z!+*26�u�P�[� �����S��¡�m�S8�Y����ָ^,�D���ja�sIŦ�u�_�|�hУ|xCgu+�a�Ȥ!(�I�6���� �kcM��q�S��.�_��r�	���+2q�����9�5n��M���|�����.t��4�oW�J���:��N�9֋wQ���=FY9����5�AAqzŗ�E���u�0��,���sYl1x���P�����I֗�v<4���owU@W��B�Y��պ��w��������Rx���.���7�t����7�:~,��p˭~���!~'[�rĺ��6u�� ���%;A���1��~e���뒜j�'[�<�z$���ɩuk~X7�k�$KGggi���{��9=R��4蘟w^���E��<)N�.�ɯ���LΆ'i w3X�Ʃ�����[xx\�:���/�C�PON�S�\R���y=d/���h 5�U����z�(���R�.�����
HHJ9��t�HI����R" "�0CJ)�w�������r�Yf��>�{?�w��
vk8TV�ʩ���t��ftx�����,�[
N�� } #��$|g�Ĭ���r�c)ly��2�أ��6=��pΔL��m�$�GS�ߋU)��i�)��T$r��[�_$c���eΐ�.��i|����[]��1��.R@g���
BɃK�j��������H�>A�;ff7F�N6�y-�7��X������4��3e���<A�l��Ѯ�� �j��f���o�G�0�_�vLW������Q�V@aK�k�T�|�ᶛ)�@.X&���N���ѡݹ� �6�v!�!�I���-�s��ܩ���k���/j����+5�k��n��Zq����;���ds3G�׽9����+���i��2��o�?
����G}گ��se��= M�o�Z��f?n�����r�o�X��;���{�����H;QX��Ύd[��}���d��pm4�3�����1�J���wʔAZ�;����n>߅<g�S��9z���W��](������8���/-����
G0�8�D�.gqH��m��U�ɰJ�P_�5j�w	�||�T����c"@h��'=!�5%ހm���7�\��b~�����X���a�V���2�QD��JǇ&د%�D�t�A��۫��fF�MY�=�j@}�e�NN��*6nF�8��1S�Ő�d�G�#��ˀ�*�T^/��F�d��<�����8 ��q��Z2���+O呕4\�����O�&������ɶ��:��� ������8:2�-�߬����<�r��9!-@J�mRq�\~B��z
S[��Ӻut�{z��V��:��ٯʘ�;٘ݘ��]{�l��d�����}R��7���B�$���R	)k C�2��8��X$��]�!�C_}��?�'6N7�*[����m�e�P���Y��՟]�����k�g�r�(�j�r��_%.��M
·�Z|��$^0ίR���Q��w�ٽc�R�ó s�����&� �͖��v�[jJ���Y��Z�����)-��T@iV�ܣ��~~Y����>r\j���s��̪�c2�e�c��2�p�n/�O�ڗ�U��M�'�Ky�*==]Q�>�	<ds���n׵��*~T	��ME�$�<j�h)-M�����2������EX��C`�S�o�$� �Fv[&<QT���"��K�<ї�	r��`��\$��f�#D��ߥ���HAV?���\�5k�5V�p�:����E���9I����v�
;���3�������p ���j�����VVV>��L(J�juO�)x-��0�^�KaqH�t$+�9n���r�=Eo�Em%F䌅"��ᴷ�UA�&��tq��#]�z�!ul��U�b1 ߿-퀘~�UBSV�)vl��Y^N�c�JI��߄e��˻�{o56������}Ƥ�[l)����rd���q�d��9q���_x��eh0������D[�1�<�]kt�ѿ��/��l����M}о0C�.���F����
ʣn��W�E���9�[#S�R����َC-i��*����&��O���%V��#JK�����ȫ�4��_���_��Ѝؾ�s����:n�~����l�J_�+Ji#��8Q�;k"&���Xx�^w|�� �o��Q��BP�Hr�c�"n~���AWW�&
��	B{8jobq�/w`}0�����dO��T·�����<<�Nl�U���5ߪ�:�;̴�M�����3��]����:��@Zh��Q9�4��d��*-��q�lj��_f��,���Ϭ����4��ci�=Gk"�u��퍾�Lo�������⌎x���3��_�>��Π� )��u������ҏ˲���� ns�ׄ��t1����-��!q��=��BQ��GGJ@d"3����C!de媡��1����~w�?�h&�&E,��G����m����M@��fM s��Ng�s�:%������ڭ�o<��ee��ml �%�� z~�6�p8"V���h@���[瞯���滈�_��r��� �pk,'�S#����\��!��k@��� xc��L��-���6P���RiiҾРl<����B��4�<匋D:�.���wp�0;��l��f��Ⱥ����EtY/��@�М��h���Ғ��������w����o�w�_A:8ˁ
�F�ffpp�����&|��ƍ�:����r�Y@'�k~�_�[�A�VIhE�];
.����us9]�~c o��q�>�)�D�
����y�)�NMz~��\d�͂o��hph*ڣZ� ���	����z�)<�eS�>=���6L\���C�@���B�I��|\j�u>ݾ�Wh��Ӛ�𒎈 Q�$�M/1� ��B2��Ǒ5���Np�|�XX=�V�k��v򆍈�������J8����щ��=qs2w�p����V1�0�]hx�[�(K�Y��ۨ�ZZx�I���P���{�k�Ѧ�R�ԥ�_o����͚��u�%5��]�h${[
3��/��J䲧&�����bh���@���S�3�:ԉT&��FfOD��C~9J�P�~��^|�D��'k�qqZ�ͫ��̓�1'7�e|hp2�&�4���(��v�m�X;���*�pKKٲZ��o�cPű�����\;��Ԋ��>(��݋�����˥�?�5E�/�+-=\-���=r7��8���I�S�d�}n�>�Wv�����1G������:�c������W���>hj�e0!�}6��8ܾWT���w8F`W(&&�4���B^'�����V�����Mfbjj��9゛��@��$��p�c���M
�QǪ�ue�D9Ą|E~ɠ�G��rn/}��g'D�u��X� �L�w����mo���|�y����.�n'J��r����*m���p.7���FȸJp�O���������C�R�um�u-?������~�#�9��{⵩�~���)"[���"B<ى癿?��zn�)Cc�X㷶 }��k��GT�����s�{����ZU���QG�����\T���W���������Yn�y�U;ق<�7[��fB�AOZf �!-���a��_+���m��X�ҫ��9���<1!�C�
¢��@ s+��su��=��'�z�^�C��Y�CW��	���o}�����ӌ���m4T��Ws*.�y�=�p62}X��<�F|�S������hDt�2�!{|m���}����4�b��|}�[n?��)��%������#�h�<��KҀ��ʨ�'O�eɱ��i�G�fEB�z�����:�"��3j�<Wu>[���)��u�G���{���z|�Jx@�}V�_���U@%�ra�k	/1���̠I��G=��8�ԅ6���w(L���`�bY�x��C��#Wl�=֊��]�A(��k�(�L�RM5��u*�_7���Aw�<��	_{��<�}~������c1��,Yv��l��4t�{���"�j��}��nB��@��2)�JE.��n|��Q�l=�4'Ue�pޘ��ࢢ[H��y�ҪkkÝ`$A����m�W�ۻ�'fm2(�͙��P��x��������OS�%��������0.�9�y��2��t�{�q.ք�q���A%[�ڎW� C�$Xp$b��,j*�{랄Ն?ܬx�I6WMF�i��LQ^�śڗ�V�g���߸���*�:�(EȌ��fE�أ�{�3������4���O=�GK�}��X�����q�8௴������^6�Y_�V�	�u �R�2.i@h5
3����7oȇ�=#o@�z7��@����:ܺ~4bk��5�T~�1��)'��|	&^�XWa^�!?u�1�;��|A ����FB&օΘb8���\t�׀E��N��nP��`�rr�$��*��� �8t�z���|���_��ڛ��_�d�=8c�A��~T(��?��wI)
��d���啕�'�k"�����k�qs��ww_IӚ��·oV?�J��_113����Ԓ>5]i1����v
���q��wu��]��w$B�p)��2`K��	�R	7�=p�cy$~�zl5��)��#^��S����j� �L�M�fb�$L��.�	4�|�;���.�XƜ%�p����Aو�L����Z���a�|��B,)�E��]�����q70������\1s�C�Û�z|ፍWpJn�;�X��������.r[=���S��W���kۼ�8g�w�`�jRX�=��/���#*w>�*p�p�`f_6��v�������.]?^B����բzI2�u��ݽK�DME5,��� / م�]�����r�;�e��L\�u�O(��@>��ө0 TV���1E~u�������dlL�Y�GX��-�\6%]`�q��$s`��L�C�B�B���k����a�����)����]�*�7��v���%� ��ϥ3[x��7e4�7���0�l�o�O�Ă9썑N0h�g�+��--x�ӧbhAҵ5����^��������g����,��ݯT
$'����%500��ev����.+�Z��s�A��N��������C�]?:�d4�p�ꜯ��QDv���Ӏ�T��}�C���#�6�(�^b�����o���vf������/��w�s�zIY(�>sG�;�e�q��q��0��׸,i�,��Xd?��'�v�*^�[I~�1l��a�[�j\ɋ����n|���Q����3�H�K�3U�[HL��5����� T�7l����F�]ֿ�{_G���#�*WR�t�` 6�`��H*"�.�<e�B�Y_�
�}
_�����Q�W���k�-E��W0L�w�@�ݱ��@�pP�k����eQ.7(�o��I�f� 1�ߙ�hVE���B�K{�zx����*yј&C�D�m9\����]�iG`��/�N�e^����S��o�oK���m� �+��4��/=��vln��O��^�z��ys��՟?[��d��=<�V�����!�!.<���|j�@>�zC����4���� ެ�N*��	IP���vc��8���cm�,|�\�R�/%2;�%�D��
E��xa�C�gYM�}Ax|�<����y�5��6�%�>3Hew‸�@���&��)	���A�;Hw�1{X��0�36q%�.�_MB�Ç��@'+~��8- �&@�>�v�UFD��I��6J�%��U5 �J�6�/_�
k &H�-����>����d�O���c�����1���. �CHx_�#��>F��11���ޤT���!145�&ڷ"�����Ąb��bw\�n�����ov0��׷���K�o�[(^��9b`jJ�8<Ħ�7��|:�w�����A��T744L:"��m��&@l6|��ر>�q�Y�H돫���f�JN���F�=��,��G4����x�m��eX�{�qY@|3��o{!_;�g��ϟ[�H��a��� K�ګ%�����rFĲE���}��\,%--_m��2'b�;�~y��'"�'�Nk��^m���22�[����\���(�3o�?�!�ӧO?�I� ��GL4��E@���j��[c�*א��L�|.k� �h��ꬻ����.��O�?�B��,�!�@�NOZ������� �Љ��dk�r8(J����Z���)�rx~{nu�W���B3ZY�!���e?������m ����(;��_��ۼ$����[��������;��8ɫ��"22o�'����G�e��'''�"'0{�<!��_�|IZ����y	S�u��f�����}���.��K]J�)���Jה��J����U1G�٣`�C|"�P�v�<!��o6��{�=�֨�O7fr��5.Q����]ܼ�LN�f��M���r7}e�����Z2&!�^oMY,��A�������6R�[i��B9զ���o��v�i.�ŞtܾlG�*B�2�f���l�?��W#�%�Qj�oi;i�`WU���Y�W�~dk����o̞K�Oe�}5�G-8�����o���̪��U#��W�"���-���"���f��ζ��}(��'(��L2x��8����@��CE�]ŷ�6~;(Ւ*Y���6A�����
���X��e'Zγ_V7L�_B��fW��o*�	�I��u%ف��ٶ��bBB�����1�~)$R$o�fV����%�Y�k���3Su�=��%��T\�rL�����M��.r�R/�'�./_b�@���ӏ�ŵ5���h":::�\9@����%���e�3�-|OĚL+�?�tR����bFōD2�k��J�Ԥ &���_iz�D� �"�<����{{��������b��{���F�&��0����VX�A�XV���8|�4�>�� �rҮON>;G~v�v��P�$Ƴ��8��d�(G_?q����~�J�Z%�n����:̡�4�/*WFӹ�����4��-K�}�?�R�w��V�`{���Tb�׶3ƌ��|",fvw�!�e��
�뻍�4���v�z�j1 �[dr2��$�7OY�q���������ڂ�&^626�y&��1�^����H��1�j��>cv^^p ,*|ိ[���Zi+i����'�[(���m��P���}u���⥦=�qq!y<GT����U9av� �DE����=����^+��2S����&6��^���k��?�����C=�Zޡ%Ξ��Ŧ�h:K�p�Q ���O�ޘoQ��41�O���N����1��
@B�8�=��U�굯���3�yP{��Fөb7T��фne��,zy	[�x_�V����,���Cž�����ag��4��
���E������\}����f����AlQ�S@��B�����=��%`@I�3GC+�Dɚ* T5��a��4�D�� H�%E�V�����%eX'�.؍~2�PiC��՝�zU������'�y������8���b�ru�`z�~N��uP��u���Ο��7U���PV���H�5 n������k��JF�4��iI�z����Du�-�������{�ӽ��kNU����g�Ƭ95��c�ۊxO�Ͻ��ُ4ܧ�%�L��˔�'#@1r~MzXc��h/����&��ft��l0�/2��ur{���66�P�I�h�q!����������w4I�LE�rrb�K+���C��/{^�l��ܳ���7x�+;/�`�~1��9G��;��L��p0������]///���F�+G0�92��n�L��C�'j�K���r��l��rx,ɠ�ig'.���V���ur+��f-����� �߱��^RAe�}��D�E�2mg�?FBt�İ?`��G�f��Ȝ�+��	ܻ�AQz3b��tb�Zة�-�)�����^a@��I����D�`�c�$f��#�.��\w�z{[�',n������ň���L�倿��'k@�F�epF��L��?|l�����J�D/A�X
,�S|(%.A^I�
Ǘ=YX���I
�E�@2��牯�]@luƚ`}�&^��q����-R@m����DDuw�"�Å�*؀�VTV>m�����5�1H�g|ʑ(Z����Tm(W1��O��@���7�t�\[#�2\*j�|�X�T�� 6�%c2�4�=�d�Iخ )��q&�@ 9Ȃ�%����/p|_�8����k;�v���4Z����j8���}��晙���j�[p�#��[���F������A]-���ל� L�ܦP��f�1��j���8ς^�o���T0f=�*�'��wTo���G�(.C6o��m���a|W4�	ɀm���"�/Q2�J��041	�"�\�΢ݱ�c��L�����v�фHe���s���J���r��T��A+�v�٥1�mG��*��P�C��nE����gS�MLL��+]x�����:coR�7�p�����BJ��r�Iti�yX��(�z�֦�4_w#�7�B��6o���'V�����/��q5i��$G)�����8X�X��"��]�o��E��R�+��苡�1gg�Y��� .��B��������W�yP��N���ǜ,1bp�����n��+$Ȅ�j��^�b_��A�Ȩ�K1�
�,W���]���_�?��ȥ���TxiCP�3	5s���jo�N4a`����tR�j������n�o��r�ջG�����WX����ZoD��� G?1�<`�:!fs`˅��}46�t�wt�	�2�����U�J0-{6���9��f�(3��k<����,O�������#���ͱ�5�N�=y�˾b{�w�9�͎�ȝ�=U�C�հ#]$�����Lv����C����1��!.�gT�*�9��t���cJ2�o:(1'ggׁS��o� "zX�e"���w;��&�JJ���Xz��EDj�W���N4Fn�s�#m��P�c�W�4P�Q�V�ܽBbbq�۴_f��W�ڄ���I#M���;C/y�]��3?��8y}}Z���{���l��8�b6�UR,��f��s�s�/7Y��a�$z�����<%%�s1n��_1�l�!��iii3��'H8�*6n���@��a��G8�_�� |�q�lj�+1�����eUlDg%�C<��Z:U���\)e�fgg�{4���|�'��Ϗ�8�8����9�
=����� ��.��c�,\���;O���9|{	�ڃ�~���� g��}Wƨ�� Ui����ss;''��^��|F���P(�+K��@I@;����m�)x俓3��}#Rk*�FՆ��f
LB9ܧ�ু�;�!nf1�}���:�_�;��G�3��uQMNZN���#���"iʭ���B2�	q�8\����+X;��\�H��[�'.�a]gQ�Iaeݸ��@��g5|��1@3���6��c�	��oqc��W���Z0�?H����^���gFL_l Z�U��	�?e�L����t��{��FB ��d?*�\�+�g&M����}����Ȩ�Q~�2I������������9���O��=I&&&�7Tc؈���P0���]y_�~q��t�c 3>-�L;��~�:\/q(DÁ�}�\���+�'Xn"����ݕҥ�/]� W���b�����{�z��*O+r�/:6)H'M��KB��h�\�u{H[M&OA���t�^�0^0��\���qo�ZEpݗ(�Q0R��緕�ݵ�3{|��XO�lDHF.ԍ-+���1��tx�;m�e�D����̽lg��<��B�C�周f���������罰�/Xۤ.���%�' ����;���8�3�Z��2̺eh:4�<���~���	� �`�Ŭ�/ވ��32RO�,"�S{{�Y<2r�>��Z�v ��Y�`���|R��h���~��KM����b�^���y���[�Iн�*��#��Ԛ�܈�+�/@����|����K+%��$tigN�/�sM�N���Ƿ�i�����l��PRr�9�=��)��˾z��eO̡t��ݽ�$Sw�ލ�Y�15�	u�� �77?pr��>�&���W��)_�C��y[U����@	%��h��+y�t͙���5#c�Ml�a�ׄ?�7tMB���E�L�+
�a�ڏs�}7qS���.//�c
N�ʔl������'n���z}�ݠx�%Wd:' ~ȶ��N��ɗ���	Ω?,����&�eБ5,lJ���ۿ��s������T����Ib�u����>��T+~�t��n�Ie��xK,�]y|�OSp��Hb-�M��,����!�͚g�9.T�Ƌ �D��*�J���-f=W�ua�'�oq�ѩ�H���"�+m����*�.�� ��{ו���N�$$%�>��)�X�|����o�ha�_�+�ƽŭ��j`Z��H$*NWK	**��;�c}gOq������/��l%�� ����V��NS3�g���v�\||2�6�a�C�E�~>��d�lAOn�z1G�,]Z������3_�xm�A����Gf�3�K�6�2�f�?D��tRWrIG'�x̉��Q�B��e��?8��0� �a���F�g<�R<[�� ������W��@��HQ�����HI!#J��7�Y���f�2�[�b����AE|��$����JET�ah�W	�ZZ��K���B�Q)�w>�w�p�z^�[c�e54Š���k�δ��*�U�Y�׻M���P�®:m�_���`�ퟲ?H
	E����FR�����Za��x?��)��nT�b�sW_zf�";u֮�������C�s\����t{��(����'AR,�h���_��\�&(\�'��6�X�pÍXF�\�ѣB�W���9:��J=)h�� A:�Y7#�<�4S<�C��q�	��~�ɴۘ���]K�țGT�����
{�� df�~k<�4��uӰz
��^�`���̳���YcG'^�*��N�OK��V��W�;�=�ܺ�=��]��F�����~�AY8v�L�eu�V�t��b�X?������T��j"�텴��$�#� V�KG��W�nk��Od�;`��m9\�n]4�>��E��)���+��Ȅ�E_>��֦���`�R+�ҥ��K���55H���Ygkhj�v�,��`���~��w(�2ɫ�E_���v���G�]�s D�&ܶ�o;���:�N�L4�������������W��$$$[G~��5P�l�鵋/5��21X��(x�E�R=.� �{y�lR<{��F��qf����K��������Y9	���_���pN��61���d}QN�%8���KI\�XU��P�_�������&y6K��z�M�)s*0�x��3Ym��7n|n,��N��;J�$����$.�V [:�����7H�}�U���m��U�"!<4��K-��Ʈ��@{���|��d�⏒R� l�r�Y|�K�r�+~t�o���@��;{@ɼ�O9�����e��Pҝ98`U|W��}Ax��
]�<��z`���Jcm$��t~Y�+-��"�P������������MQ���{,�y��G�����zO�Y�� ;��2 �X���%٘J��Q���`C'�__�uX��++W��wh��W=L{��q��&$S���<���V��I���oQ����C1�W���!��B�8&�7Z�X�dX�Ym1�gm��nք�� ?�+PR�x�:|��3YR�?v��C�]cF��`���-
/)OꉋdNz͟��jԣ(�u��;f��r �9@����ń��_iyU��J�饫k������!9@@,���X���n������vihk�͍�<����ʥ��u:�W �B���A�v�| p�±��E3����������7�U" �}a�� ѫ�����䃓�����+������a��0�%{=%ʛ7��`�/�5T����j���������8v�ŀ���"�M�"��KZ�<��g����Â�>��B�v��	}~�l�\kYѶ�B��}n����?���=޲:�a>��R0�ϟ���Um=��M+��Y�����2�eq���ەy�����ʼ=��Pah��¶��V����}�k��]C�n��8����s{�푝Q8"Q�y�ƾ�g��
['������e�����:���6���mV�苛A$r��:������%��~UD�VL����7��2�˃���|�(~�宀@��a�r�N������Ώ��j�G5����SFG�����|�C��䡀��d����R^Yi���7�y;E�ϸO�m�A��l��V��ss��cRV.�Ý�@���v�����dg�t��\O6!@�A�@M�1�0��_4�b�I���w;�Đ~?��|����)=c���5�^ˇ	�d�����de��釣0�˾R, c�å��q���|��er%�� ��[���5��@9�h���0�E,���B��D`ܾm؎��3J��/���(��ؠL�.v�<�V[~�$���l7�ᗗ7��T��¤���»��λ>��6NK�!!=K�Up2�s�=�J�C2缓@��2%E�C���K���tY��=��ϊl�gGFn	ܻ礮J�Dh�66���\��o|,�L`|Ni���M�3;�--��,����n�� e�d*��,7��Ȟ���w޿� ��4u�����\����x�5��#T !+� �U/
�#H"�����"��S����_.�D^=}%�����i�K����o1���n�,�͗��D 9�ܻ�q�l�:q�OF֧��t$Fs��G��R,�of\$��Sū����c��vKq�i*tb=�y�,
|�L��qXz�EwOD������ݖ�����14M��zv�'	��*G�/�k3�/��˓_�lV�hV��द��n|�ՃV����`��=�BB�Əy�n���Btw��9�E�l�������;����ik��?j$����iȒ�Y;�4��2M�}89qvqu��k���;�mii�GB����$�ܿ�0��[��0`���������]3�_:B̨j�܄X�c�w$UY)��e^h\Q��W�U�V#�^���1|b���B�1����z��8��A��L䘧>�a��qWy(dݚ*�6-,چ�f��/FJ'Uw��#�W�Q�0^��ѭ08l�f7+fW�r����9�g���V)�90�]���g�߈Y�&B�v�{�=�_�=���@iARN��v��d�C�/%�3��!�3�3���3��ȯu��=ր�b��9O_AYY�ڬ+ckd�UU�${���d��NW�x{��|F��CB�*V8~�mI�g���ҠJ���ߊ�c�uDȢۨ�x���?��G	�B���ܟ>}
[Y�I�'�o_Ѯ�=,��ԜxƇ�A`��*�Y�oVU��;s|L|��oJ�&�J�n���[�� %{z�r%�_��4#�����H#��>%��!����"6(��N�~�g#�R����sں'Wg|�7/�j3�	��"��Ӝ�6'�i~�k����Q5�h<��Ƶ���(_�;�R�S�=��n�7-��C�&%�"(G��z:/���`6�!bsp����vCN"K�WIIv��{���T+^P�-��z_��%�ͬ��I\�!wrr2�ћ�����������;�Vܷ�����4��,\]�gV�Rԯ<}:��CM���=�xv%�sV�~Z�����&!��R�Y�D!�g�!ߐ��'i��-^lD_t�n�% Ǘr,1֊��}�Z���29xb]����"�}�h�'���0���^�DR�g���.�$`�|�5
�/C��ҹ\jP�#-1��sƓ������	�C	.�̞��0{X=+��I�w�@V��T�Kr(�ݒV��[u%dEo��j���<*ݡVxT�r�+�\�f�yՀC�^YՌ��z����uq��lZV�� ?�8���}3�?�GnLP�Lk��$b�{ٿ\Z��"U�,�	~��T3��02>�dS[[��X[������
X^�@m �h�s��D]�+���ѥn�u3A�
3_�i*��ttwEF�{�X�=��[��������=@��҇�ݾghMO�"nʸ��C������Wk��B��	Jx���������ʗB�u�K4akDXV�k;o�-���r�@��� ��_V�p�C}���+�4
��hۧx
肍2�a����wb�������o5N�)��{P�s}[<c�խ�81i`�Y.�i��>Vb�W�.���ey.��c��l;ٯ�f�{o[�t�4ɔNm���k������Q �3W�b���+���0UY������'��rSӁ���4�Xʚ���R����FFJ%<�L�D�/�d`�g]b
&O�KF8�>A7� �4��j\��������A����i�XV����ˬ 7q8;^��U��<�]�#Q���]�@I�*��_n�K5@!96����y�	&�Wl�t�Z<-f�]׾�r;U��:.����t��J�*�m��w�uω]�(6"J��QjU%�qo${
�Ԅ�ˍ���?z�J�-X�<8Рk$-t&\��on;B��.k�(����bV6�B���}ڬ�:WW3W�>�UE�;{6Oڂ���/�Q��N���n����;z��k>�0<<�:�h%պ;����pGFCI.("��}���IIX�9���}q.M��<�Ŋ�#b��.����?����J��ޤ[�*Z1Q]�c�M)Zg,ū���J2J���i��G;��mJ"i�#?�j��t��Y���9������)��s\/�n}=�8��ס*'��u�0F�z������0t�ڶ���G�c��ԗ��4�My��Z0a��$�b�xl��ݿ�a�sz-��K3pS�q��0�y���VwOr�c@��b ޠڎ[>S��C�ʎS����nS�323?KE��{V��0�S|:�`8�Խ��OmGo"p&��;�C����16y�L����&�A�'�[�r�I_��l`����5;�+�!
C�6�^�=���--rᕌ.��Qsg� �̪nD+��YS'q�8T�q��q8�89���.���|�n�Rm('���/��\E��hM'u���7���Pj� %[��6e� iWP%��)�� ��ZE��V�5�?,7��U/r��+(�/�+V�ӽ��`a%�$�i��A�\�S��m/��^;h�.(�ԁ����`A���++N���j���΂[�:k�v4�*�������7+�����N�ґR��R�kk$�M �rr^��H?&*{Eܙ�hP�}v�@4+���pI��૥Џ�� �g�x���G�$����rk�,0�ʟ�Kp�Nj|ߣ��yݷ�')\׀�/�<AR�[�@3{o (�PK�M+o�:�P��@Tl<EL(UtA�������ط岏>;r�@��p[����O+�a�M̝��:�v���2�A���EL��b����t�$�k�&?�l�a���Ɂ����g�'�ퟞݿ�
_oS�q�I���V�K6�J�������ihb�9[�t]R���?��3m��'��ܦ��� 	�H(�ʬ�<����N4bo�L�)T�����s!j��KZ�Ǐ�����U�,�uZ'���#& �r�~������A ����zx�3����jb� 0�WK+�g��I$�E��[׊c�@Nלﻌ�c��k�����h o._�g�e7��Ł[Yp����ae����C A��MhI��C�.|"�!���y\j�e?�N�qt�e^m��0�<E�;��������v���.��!�.z9���^��UnS2��U++ī��̀~n�ߚ���؎1�vVK�K;VSu��v3��Ŋ������SF����
)��Z\]j�]S���olr�G=���~ʰsM�i/���P��%z�Κ�L��[R��sD� �ӵ���'&��3y6�߻�V���Z��ߜUmH��MM3o�֑=�6;-�<�C�Aӥ��B~B�=Q�C��Pyդ0�j��֢�#W :A7R?��i����$]Y��Qv�h��Ika{3�OF��rL��'������k2&Kk�)�C�|�޿�32R�1*W@׽c!ë&W��6��W���Û�V���.��B���N�t���c� ���ǂ�穚͛S9�f�\���w���.��|�?�=����<���qu�<姶sj�*T���2Α�T���4�v!./_b�xA�����{KIX��h��D�Y���J	�H��o��b�],Ñ444� *�wi�>pK�^q�cT�O��v�X��A��@��N�hc�}<�vY���ݘx= ��Y��{ ����.���]a��F)���1	�0N�S� D��@�➗v㤡��B�׋�q��Ƶ���x�7m�Y�E�%���&�&���4A����k\ޤ��ש�m�p��Z�u�Zq��oR?�cOp0���>����`zӆ�����/nU�B3A~r�5�i�a㮸V߾�>�Sɝ$s�g��4!}�)��fT1���~�5��; J����Y�M�@l�v���7UG��+a���c�7-���===��9��K;~~�u:��s壗�22��Q� ��_��5�+.�堦�''h~���������f�2L���r ���d�'����>�9���Y<{z�DHx�g|��ѫ7J�z��GG6վ�.�39	�_�`V..�]]][�-v���?
��W���m:>����X��e�N��{0/--E)[�
���l4��0���[���+J:*�����%��@Z�<C3j��H{��=u@�Q��U��+�ŝ��Q/,�<z��m8f-5�����6�RX���=%���o�A��R�n�{{���Đ����6���k��{��~�3I$"��כ*Ƒ�MĐ��#�g��F����A��u�razz���;t����V�Zy�� ���\M�U�|O�$�`x���}a��o22n����Z��~H(�|��&�g/_��^�M�:�h5S�e)�(V�v[6n�*����H��<T������Y&��5��31���k��;S/��Öxl�5p�_ǌ27���(n��J�9S�������%��^�ȽzuR��Ow+��4t�6�Yo�Yqg���"��C{Efzƴw�d��qCU!Ƈ�#���O����D�e�idf�cN%)�Lw�e�է@K��x��O�����<�a�����^�GtmR�>�z^{���4Q8&23憆a#�+H�� �{=������5�7k�[&�<ʳ���pw�M���Qp�v_�l�b�β��i�����Ѓ�\xY���@A�W
^h"��2z��{PTS��DY�?���vݓѳY���Q�m-XV�D�'4�_���������Gf��Hߕm�Ev˱m=N|pq����J���9 ��~������T]9*9����`!s�6]����{��+�]�ٻ�k�t*��Fp�s+(t�jd�h�A�Վ)J05�+�S�9}A]�պv쳾�)�NV�ƃ���3��GȺ7)P�[/��w���q4]�lf� ���K�D�Lc�{��O��UçOm�qqq���$(@8NN�o����}q�~ci�)"%e�����<C~:~�f� ��z[+H��L$����B2���/�N���?���3Ԍ�zzAW��q�,"?��:r¯NO�"�q�v�r�Ɯzff�""#gݛt�F����J�~���Ҍ6�L�[#��Q���.�6	==}GGG�Kr%��K+ ��[u����f�rz�Ҕj��ݔ���M�]Y�����|�yV�XI�B���n��u��u�ؔ��
�>�?���v5Rt=PHJ.��]�,L�9��_��\�+]W�&�O�{�]�����32��I��4Y��/����Ĩ윜���N�^m�/q1ۻ����ѧ�Jf���xSt���y����ۮ��{M>��3ss@��9l?x]9��͍X;O&�iv���v��h:�x*����B��!���#�Yɱ���cdfo�압d{&!�ӡc�8f��]����?y��u�������k���m�Jԧ)����"��yw�<�{�8��k����w�ֲFuR���DH�1T��������R�lT���N����C��f��X�ʾ�j5�,k���2�@�H�M�W�ډ�-d�z��Ӣ�y�g�|��]8��Iĵ;��P�Sa��sqi�Jk�a��]�W��u��JZҋt�9՜�����@VX�$�"�e��E""�&m����h�[�##���34�Ty��	4�y`}M4\H�uE����n��!D�m߾񇇇�㆗�nl0��i6؏P~Q�fl��I�+��,�ֶ�ʦ��#**�{,�=�Z'��ח���W����o������IIt��鮸ջ��θq�Dqё�M�s�����*߻)3Ʊ峩p+~:��	u�����i����ӫB�Sc^�.v�o��B�����t�N%�RYt���+�q��V%=ŠKoP�θ!��<)9S4�=�����	f��.Q�7����;Da\k��<F��9m���k[;�Sn�pYG`p��Ke��,%V�d9�R��z�<����afe�z9=�t$����:�LŮ��(�(b��Q�BaΠh~�26-��n� D3F�oA��hu��F�-���G���?UTl)>��2�@���6p9�Q#f��]�f���_����J\Gj�A������:��ƥ���
��n���xE��Ot����I��h��Z��@����ß
m����*3�'���K��p&u�yh��Y�vfvvB}���%3��8���f�̄X8�>?�^��e/�B�h	T�"�V�p�����dy�������ȗ�Vh�%�m�8��4�2�}�[ƽ��o_U��<��0�Հ�
����+(�a�O#��a�H@O�үyN�&d��u���l>�\'�@��\S5Ӵ�X�fSh�0�sM���2��ۣȾ��������O��^B��㝔i`�������@����Дd�ۢHeKK���M:��_:p����B�f�i�^�����]^P��/)2_:Z8e�7X�GEF�y�p�]$E��R���b1E˔�����宮0ꪢ����Ծ��q�v�]6�©�E�S����_嫪���nlZ�Ԗ��p%Fn~ 0s-�N�?'�ᄜ�Ǵ�!�D��jо�����.|�Lj|mo
���TM�6��k��`l�K�T�M<����̫[Zz��	�#��Xht7��e����.������h���+�&<�ƻ,��0�QvAA��w������v�a=�e��C"��W3M���H��j�{�,[[���"c��wɑ��& �!��Sh��$-7n����ù�1���?B�Fk�C���AoRp����^9�dB3�MOrt��̘��������}�|�٭�͍����Y�/|^�u�.��m�>ZT����QP(���uJ�2�K�HRSD��H�s8���q�@=[��v����!��!��v�*����!�%������V���*�luo �-��*�{�b��GoC���keP�	*	�!~l�1��������k�T��_ut�薹)f�,5L{{yED5��R����%I��dL�G䨓۪���2cC͐-���b�/�М��L=�A�o����}����`��z�TQ�nұ����m��TxhR�DP_b�ld��yH�f�)tp��>���E#ߍ��ǌ�pӥ孺D����	���}�c٪�5i������5�K.�rbi���S.�(	��)��ʏ��i���3j_dӵtg����A�+���5+/g��XR����9�Eu�v�H��`� �&�"eÜ���2ܟ"		y���C�UL�<h|��.��5�ς�p�8��%��Eb��]]���yGvk�������W65E��Z��@C��x�uXՌ絘��J��Ķ�k:H�����WJp���d���o
�N)��wG�A�:0Ӕ�q	�k�<oE�8�PS�n�Ȃ� =��^�c:a5F�o�����IRdZ{Kg�!���l�ۋ�w�*��T�<b}u��@�cx�ו������e`,�h"i�	a`�;(��J�:���jE��$����n�<�n(..�QgN�^��_�qKU_TNNď�ؑ����XJGw�D�=��s�	k��q)�������n���F��9>(Ywq�����KK�����v�=���O,w��ma���&($��Pཐ*��t�D�ľ+�8V�oZ���n�ݓ^]��y��q�8B��C���ʶ�ë1�J���@��W�w{�(��|�^�+si��C1����q����\�ӥл�Vj\
��-l�׾>���̸���5�%�G��?��h�Ԏ���5O��4o�(��:	�N2�\N{�A��G�-v��.�ywy��P *I�����L�����+M�U��my������������:Vu��K����D�#�iO��R$�g|�$Pi'��M��63<<#��Ɠ�0	�<~^��?E8Y�<w��2�~t�bP̃:�j��o��>]�@/����~��S�N��P���J�k�)xv���z�>?��.�\c��O��"�����gΠ���
�#��P�N�������&�4�ʉ�B�?���93��a�]�%�u
ݦ�-���χF��ǵ�c��qо�+�Zwň������Ԑa4��O�@lԍ���Q*����y4��_x��Э�;=���׾Z���A!*)���}*@ղ�\L������b�(ik�/����7=mű�S��T@HDTU��X:0�Dx}����9��l���^��J�>����� )�L�+Ƿ�:wr�����Ӄݵ�،��&ip�M�Y�$%��z�1)ƥ ǵ��������3�������;��շ=�Z�w��oy�=HS�V�ֻ�d!%��0���c%��\�R��7X����b�͞.i���)td�P�n_�����@���N�9�C%L��6aj�3P��
q�9��T�����
y��~���>�+��<>Й���p���ϘO�Q�XZwvb��ʝM>T+�fP�߿o�D䙧!Cڠ~��=-��n�y�r�O��.2�� C�*�ƜN7Goo��ǅ=�#�ӣ�����I����k2U�b_eJEF�t�����3SVM8u��;hX�I>�]|�=!B��A.�%-#!a|QRr����_�
"`.!��zt����Ǻf���?�1�y�(�9��^�(>����N�f�d�K�+)���-����ND��:0�
|,wo]��g�~r[���,� �}��h8�p�Jf��Q�-���+WWe�ˠ�A�vL�զ��,�J�u��� ��}�wո���*w���?>��=h����5!�By%H���{�%3��������OdZ"��D G�-BH�-�i[cFM��V��hȡ�;8 �'wF?'ٽ�,h_t�D�,IV=#���;�^H�B�����zs�b�I�3Ow� dE��3��kj)v��0�Z#8�P<Է@�X�XIPq$��R��Ή�8�sR�}�k�c*�6�����ts�"��+�'CyZ�t�t��(X��E���{��ɠ�U턜����ǵs1j��]����nn�S_	�G�g񀘥m�=#--lp��|��Y�n��(�6�=�-�,��xH�ع���T;ji+�u���� -\\��	������TH9:�	[�D &  ���N(h�?�42�{B|9�.JJ�_f3D�4;c)9W���wr�e�y�Z�Y���|򭎯���U#@Xٞ�w�a��z�)��2��V9�F�CfC�#1�����Z�G���g#mH44�����/����g��~ީ���f��������|Fژ������\��"p:�[������K��N{�`��f��@���}���|�[���I��/N&�P;|k�r���,�\��9�b��	���b�7W��;������Ā��w>�j�!? �.�gܨ��G>�b4��㡆��e�s�WRh�|�zն?�MZp�R$a�_��6U��{#kG>�ZvH$Yt�X��p���0A���/#5>��s��<��C�x����}8���p�������Ǹ�r�UH�RL�`��`�@N��3�����^Q
mJ���k*����g�[�Hķ�A@��ܑ��.z��|	��<{.�055��	���{\U�q�n?sb��Y�p��t�0>|��<�� ��dG���S�Y��
1��T�֛�6���jrh�۲��4ҧT�9w�'����;�*Dޢ������L�$��ȸ�$�kp��S!ޓ��5f��x�cr-u%~:����@�@�Ix�@M�\�u�2ի@�o�z��ғQRާ�uK�����Yg./�e+��%M˸�Cw䋮����)4��ʛ��S�l��gTԽ��١�ˀ��/��DLWpZ������ϘؠbX!а�� 4���C	�̞���`T����^Z���qq��L���ꠅ������?�Ro�Z��$z<g���I�9Z�G���4:\�b�
t)Q����"�3��=�������̖w�I��X��> �K�|��E8~���?F	������yJdh;��
_�������^�����fN��O#��{ ��������W_:����n���E��x�>���ˠ�{��MV��I+^-�J��m�6Z��<M��ށ�k�|�2��"����N��ڰ:�#l:�<Iz9x�[VI_x����u�7�o�bt,ʥ�ߠP7}���JJ�:�1HNFv2Z߄��K��������)�%%�15�y^6��^0ۗ�r�W{~��u�O�ࣖͰ�C�F@@>� U���l�gd̅M(Zk'NA8x�,���+�Ag+���RR�5R8�&�Fȓ�LFQ����i �Ϋ,rd�O'�?4wݗ��휡wʎ�����o��g<�G���I�Aֶ�AV�ʉ�@Ĉ��B�d����M��>�:����k3��I6Y��H-o�9�=Ar8��[[<)��8p�������x{�֗���&_���TR����D\A��ý�ۀ߻�x;��w�:���_Y�"Ѐ��)죦�(͢"���&���dH��
�4'Y�Fn4�'%=&���L�w�SU���zxuk��RU��A��7�_�(�1D�0%G�%V��4���
�:/�&R�`�7T�|Ñ/ܙ�l�����Z"��=�H�P�C����PS���ʅ̂�@l�u�l'�F�?����Ύ��;WMm�~����7�V䑙(�������f�,ll���A�
�M��KemoO�S�����3F���e�E��7��2���g��k�c�SH*b���k�dq�p�AS�C�DC��A���|_�6E ږ�{khh�$KJfA������嫠�=:�딀���������P�J>#4��2��v?��RzҤ�$Ǭ��%���!��R��A����a�1�q)���#����*#�B~�1�O%Y�/���}W���z>���Qndf��lBl�=�c�0aɌ~�3ʋd�+��Vp	|�d��1�E��EQ�#����ݑ̐�������g���`�"�d\������{.,�(�Ʀ���!�΄�9��'�@�����f)}�;M|!�ijn���ε�y�bi)İ�5G�wvB��YOt5*�լ,�������2�cE*�yt)��D�_���;�� [�����r܉<z����-H/4C������=�ݨ�r�ڹ��%O$��;фߘ�j�Q6��:p�|�(mB��tyX�[Ф���_�@x���X��_U��vw�`R�m�����0_�4�5i(�£�����?��`�j��ꭙޤ{��,ͧ��˹Is!j���m�|8��n3�Iw��}ĺھ<���O��śĬ�Ak�x#��ۮ�e�9p���v�+:S�\� ��f)Z=~�\3>���/����WKK�����鞒1�3�y�s);�G�uu�S��k(�b��W �ݾ��r*gPl����en[e*�x��>�T����uM��HuUCK,S���;8s��x�wq�!;p�u�%,�"�@��/�ފ������� 6^�dMB#힘&Ĳ7���}�������NJ���P�!�?�}�t3�w�y��Ś�?�fe-�~�al�j;d��v/f�	��i���2�C�P�����kFFС������p������g��0�(�|�@tpb���f�3��n����(��(P��E�D<ˮ�P�9�{G��`��w�''a�koݴ�? '��G"wTe�u$�߸
�ii���G�y<3o�%�K���HNLIq^(w�r;��I��#�d~�
��׻�LӲﴙu�N������K����7O��4�)��}T��� �Ȕy��
��-j�A���!bCF7��no�nz�ה�`�X^Ǯ�Ft��\�Q�Z�?V���Gll�ۓA�EH����X(i&%���WcV����b����;�8Bŀ��F� ���hfU�m��/6�li�C0&�QG�Ë���(()Ü�Tg�]&�`!�� ��$ ��J�(���,L��n�2IN %�O�rp�M�F��@=6�.�=ͳ�[\��x����d�\n.*��(:g�_�!�M[,Mh���$�>�?���0�D����L:S�������@�a���-b<.~=�pff����1qzA�>~��Θ����c)�	+,v���t����~ĸ�q�SS�C��/(�eQ�Aw��	��Բ�g�y|�Y�d��=��[8��u}���97��>k1WPXh]喾���M>%o�J���㒕�M�Ѱ��C*����	�+1�y��H}��kd��o+�"�"6�җ�m�&�|Gp�mk�2k?x���y��������j����:�&MM�zHr!4
�©�e�>fP<��>7���k�;��iďZ�-(|BE������O��A�.���es{���a��_�U_�FSrLnYߠb/1.5�8���6����v�?Њ���aVt'g���
�.��Uo�z��Xw�Iev�RU�����}B3B�����a�be�* k�i�§=�
��v���B�����5UvD�I��.@��u�Ɯ�_���W���w4E���US]v��+t����ܿ�}��A�mȰ�En��Puu���I|�������A����w������GC�H,����rPKqD�0f��bb�芖TϢ#�Y-�\ǔ����o�B�����k��ލ��O���_&�B9j|�+rm�#ǋ�B�M�feл�|(����6�כ��>�Xp���P���\\s��U���)�n����3@6��A	�.�Rj$��6�EI����Z�rn�|a�����A#RN`$n�N��5t�l�m���7X�TE�ƺo�zV����C��&N�h^�Frh�*����樽�G��32X��O"����o������iۉ���r�;�<��J�h!:��u,�MLxI�����wd�����[cu�^��W8��z)Y����Er��=�T.�et@Gm?tG�!�\8fd��rÓ�kHj�-_Q(�G`{�a���7��  ��}�'<��Pp�O��S���^���4�N��� ��5.�����\\o*��Z��������e:�����W�R�����Ç�;�z�w㔄-~�����i���~v;��ú����C�ml�S��F��2q�f�b����HScy���z��]���Ϊ��r��jnO�P�|�YD9�$!$�>>.�םb�C�V}�Z����"��+"%Ek+�B,q��^�^^�qj��n��G��bT����Մ#�C�����G`��s��(od�C&Q#��~��~��� T�k��jb�&H��:��#"�kv5x8���J3ā��fmӔ�J��ZJ�T��~	)G��b�w������������o֣߮�z�w7�e+�~���8�5`�|��\��
����j�h�0��B]�����}z�w�L hZ91�yLI�C����c��b��g����[�u5�[�������<Y��� ד�1�
��LDD4l�<x���}�4`c�l����-N>�����I���'�踴��-s<},��?��r�L~�X��]�]�U�T�8�v�;o�J�*�Ƭ��x����l��e���=�������.7��"�ւZ��j�i�[" .c}��-<f��[&ER�W�H4]W(�.���:�r�����3XT-4�tlE�.�M	��n��ncن�5O��޺իF� ��iZ�Ĺ������ݿ�Ƀ�(��͝�ۿ��#>$|1�^nF]*�k`�ƋXR���y��b�j̔���[�z�|��Q�Yx��;-^P����݇�'�^�Q�����]pR�?��߷n��i��W�������=�r����ǜ���A�{$��Y�6�p�-'U)�\����|��Nt�b2���[���Z[K������
�¢�}i�wJ�W�t��N�a�� ��H�d�Ι����ˋM�L��]8�T��֞��w�V���_κ`Fƻi�)�Z��+C̕��ۀ0��d��!��-.~�p�Q/�gmv�nG��V�IB���&�,��HYA:�uٻ��O���?��ʏ�md��\&H�ƜN)���6j��u���mo�0,���E">ߣ�"-��AG�1�F�fcnF��K������z� u�4-^-�AR��Cy�N��^o [11�q���b?�S=4�<`��e�����_�3t�:W*wn�'���g�R˰ B�Ѣ�/�%?	����B����7�}tG]\�>;<�_�|������:5�y�H_;�. ���"eGX!x6���ȕ*"�u%�	����@Ha\��8��]:3U@w�G��o�z�|+���9֥"�u$	�]~�ʝ�V��w�!�67#7}J�:1�A�L��"W_
��=ٔ�7�{�\�9�'`?��!4���z��t��?_Ҷ���iQqP	@�ٙ�C	�=�fzI��.��B��<�L��[��R���T`�w���(���xRcVU��f\z�z���T�����n��\?]c�S+�sH)�ܰ����Tb�)W_��g����q.A��W.��0.�]qI�E�b懲�u(F��ȗ�CM7��wPr}u����e��G V�)5�}8�����!U ��LLL R�f?q~���=s]?V"��,q��QE�$�O�ax�K�=<҈Jau�� `��p��טG�G�v��z�;Y'k�?C
HjŎl�D�IE3nŋg�6;����=��SH3h-�A�Mդ��%BSU>Ħj�?�0i(���#٫���z�%L����3^
zƿx�IU�I����1�Rv�oA+�)�CZAs�zA�n��6��Ӹk-71s��QiJ9̂z��knV��;T��c��qmU�(�KJJ
+l>G�@g�|����{ﹰDs�+��{\a�o��� �#�@;�T6�\-3��>,n1b�����i�; ��JM� �á#):��e�ML~:y�g���i��
�5f��^��)w6E ��:6/D:u��uȻмoc9)aq7a~N�XY����)�WS�9N���5�2bc#�Ԇ��5A�)?�kG���m�t�e;�θ����d�!��(���s�:���'F1��:x����zo�]6�8�3"MGW��#`3��F]������7�$/������eƤ�e Es�����edd�Û���g�G�G�����''lϦ�"�oo t���!8�"K��b�H�y��T��IPP��P�I�w�.��	��h��ѱ�/�Ņ�+��=;ğ �,x~�C�@5���䤗R����8Pz�S��[���E.�RѴ�������s����ɂ�[U^]����gV�=�!������^o�˟#>'v �{�4��))(>��(G-	⭪z�ܰ�v����n��	7�9Jw7�f���o�9V~'W-��F���*�<uy����!-�+-��c���Gm��+)$���Y�l�V�w��v}���gc]�yA������{{�u>�ƈ��<��:*ѫ�#�J[�������"��DЖ'j��e�+��v�mjw��cɉP��	.4ꥸ��pVK�b<�U'b��S
�P��?;o�k'���OACy�� �Ӫ�o���"�lR~=�~hXj��N!i��a]�q��<t5W?hߏIp�gc�}����*eoo?��؜��Ԯ3��!����wHbk;g���2��5����Ejdd�X��F�c���+�-��Ⱪ"� ,v������� �g��tt��Ș_G7�Ck��qn!��)Q~z���Zn�g�9�ɖ���"s��&�*�?47�Z���{v��9,��X�*�WJV��PR�Vq4�E94�9՜�6�{5&��n_�3��~�LO}Z��O\:���{�g�`�C����P�����6��ه|al3�?�^������I������3�;�)�(()_k^C�4�
��*_��OL<���%·r��=�"	D���#Vټ5O��ʘW�ZW�X	`fUU�P�&4K���i�%�E��S�0��s�P�0��:|�L�KK1�9�L,,��by&Tj1.ė��"�d�/�dx)�/�5`�O�/��w�/F
�C�q�_�|��]�u��]H��DT�;xQ`P��T�%��֭4-��Pg�|�0R�2�#:�%��Ӵ�!���I��@�P�,�<9� ������*�O`����b_'�E�b�v�׳��A���k��px��Wcb��d�#��lWUF�6���������>���t�aZ���@A*#�3�}7t��j@)�)��'i�XIz>S3y������1|9�F������� �Jfx��|	D�����*_�>:���h!�j�ܜ������H_�]��;	hq#?o���j��U�N��ʙ���^~�����m�}���E��^����m�
��*�q|���'�����!�&�4����Ҩ�K@��D��ԄԶ�V��.a.��А�4�&]YY��� �A�����z�/	y�K	=�w�B`\8o8*ιIS�TŠ��h9��I�b`r

���!ó@0��rCS��n�9�[ނ���[��B����wO{DV�f��q�]�5DZ�mO��������?KY�	y}��#�r�p���z�mH �����ԤW��VGˀm��8U�s43颰{�K�<���%Yu2%�6+�)�}�FKt��d4|-S����y�����o����^TZt'�$	�R�R��~����^���INj�,W��I:�k��������J��9www�t��[\�1��I�w���\޴�����
AK�5���΀G%�K��|�]j���'c�܉�׫9�4��1~�2�?�91'/n]�|��ɍ͓�c�"��~�iB�Z*|pMsꚟOFbgf���ř��Hl����ǜ@�zhF�|��O�����~I��]�g��x�|`p��]|d$�ڦ*��2��ݫ��@a&�Z��y�;��a��KF�j===�H�9��"��T���'dn[;A��G��Sw=iVx�""$.ŧ��G�6�q�{� �ԩ����JB��7�*ӳ��z@*|i���7�O���p�E-M\
�[��p����������U�5����_ye��VH��[X{�J����oət����\��\̠J��~���4��Ԥz���t\���Z�T�5Q��`E�\9�I�B�+��)��Pq���
��	�B�y��k����&8���'��_��߿�A�W07��eb��/7��e��R��1�DR^F�Z��Kr����/����i?��5�ξR?�"���P52��?�-���p�����!K�9����|��cH�6�
G��pr�'i��Q-�����s���݄uP��=���������J�*�O����55A1�0�����-Z�(�*pЂ�F�}>�b/7בmaa!^�}�s[�P�R󽳲���1�.UO��m��Gf<pB99I��x�4Q���� ���̀�u9�h'��Q�^��_�NiX"3:�����R겙)�޹R�l,w��/]^4��u��(��Y��i&>�ٱ���T��+�
�=���n���_���u��-��ݣ<"r�:������DԤ��qR��G��ח�f���ۖ��A�"��$b��������C�Q��{�0��r�aQ�����.�^�������M���%�[�hh�ɠH;��UMMןS_�"	#ׄ�.(4���75��Y�7(�צ-gfa�n�w_�}F���
��o����Jv/.���BU?�tZ�`��SDCM�p	�J��#�?��wB�w���L
�<|IuKU�re�枸��8�Gd�ڽ	xR�,�BY&4����Gh���7|��'���z����Y��C;'� �	h�+ ���J�=,���>=vL
���I�h����Es|����axw^�Ź�KEh ��&��""�X���(Ɋ��hi+,L��x>�5+��15�:�H��4���̴eZ�(�K%Իܡ���v{qw ��(���%����xH8}Rx~��b�w$[=���cڹ��8��x���u��e:-29�	�O�D�`.��Gr�F�<���C����v	�a>�ԏ8�ډ[�����m�0�\,q��)w?��Y=}J�P��:ڧ׵��q���Ʊɘ�Ɣe�aj�Dj��-���v�����^���t��%c����2˲-SSc���R�V�R�/q�{{1:#&FR���.���Ѥ�{ۦꝲ#,D��3w�Ծ��§�/��aM��^�鬟K�
�`h!��b��O�́���+�3���C˪9[��s8if��j�f�[�I�^�$��F���NN�ߪ�{`�o������ʱq q�J���{�eDR6.&�Q9J��M`[n0.[Xx\���_>�wH��M�&D�_��7�,��^GF~Ө_PzX;����S���eR"5�st$ ��\[Zbj���/�Ё�v��B+�C�KJ�e���mk�n�˻�������Qq\�_-�k⚰�?&���5i�|.Vd�5c]�=^�P����)�J��?��Kّ��?�r\�d�2��!���κqG��v������w@N����F�©�?��d�Ƭ�N��X���N�Q��a��}x��a=�b����3�G8� $�Z��{���,��o�+�d�jM41]U_���6E8B���X(h���
!�����;��jtu-2��d۷�\.(��Pc6\32r[�]3�H���b]hi�!M\�����&�����y��e8'�W���[�j���Q�6]��Vdƃ�a,�4-�����E�t����Z1�>mr9��Z`|�W��Z=���6��a�ݽ�Vʹ�v�c
^JfXS�Q��G�jk'����'���������k�	!�m�z�G����|�����K4G���@@�-�gfޤ��-�<�Icg��.u�پ:H7KqSJ����	l�ņSS? ��'��y�Ȗ1�ħ�
M���Q�,��AZ�w*Ãc�!.������1W::�	��4�[�ir���5�u�NsH�҆��e�)��߳󭕪ܚN��Q�w&r�=�)���Ż�S.��g3�RvR��7�W����UMlC��R�a	_�޹ YcN��<�:�>>��
����Y�|�I����c��{���C��/��r��l��){�n�������JJ�s@���=�i,���!����wh�WU1pr�yvK�b�l͞(�b4c�9�m,A)񇠤�Sb���=:�����L��_�aۆ���!mxl��Q�,�ٟo�ko7дC�)u��q�uSoD_�\��A�����L�Z��K�G��Ӥ�3��͞8i�{mp�3��!���.����i�FC�߭���GЛ����	SP-̾NL��`�Y[�����S�%γ�i,�P�BLX�Ga�E,�g��<a�;Q��Kz7j�n
����v&�5��>���'r�Jڏ4d�G��;+���������;��Y�0�ͅ�l��.e�� �S4�_��ABs����=�C�$G��j�R��c]��mn��"Ɖ��?ؒ�1k�s���dT�҇��AXFW�w\jU�� �=ʼ.�B�!���)v�3O�wS�R	���4u���!���~�H���F�;�/�-�fҁz:�l�$��eirg�_ɺ�0�黹��E"�1�++�"o�^6)6���q�2�Ihw��K�Z6�o
\��Ov__��Gk>�oA��TP�����q|�"�t9��֖��i^���d�d �
�9?CNFF�ɂ����yf�5�Y2���v�-����
��Qp��%��]���=%K���<$P��"��mP'�}� o[�2'כ�Q<lJ��@�k+�c#U��Q����}����S[��.�9�韭G�B����dZ���{]E{ ƭc]M���2�1����Ɯ){+��$�p��Υ�]sK�g�>M�|��b7�r�Z{6�����,��ޕj�+k0{&�HT�%nS��[dbh�����{5�ܾ]H�|� Hc�		�΀�G
G  R�@�x�3	��o<P��Ⱥ[$�,�A�km�"�8�=�����u
�F��+�f>O�f��_�Τ+Z�E���qY����Z,�mjty�**��2�Xo��o �$i��V�q��4���ͅC����i�#v��@d������M���sjc<��m�TP M�r�2���W}~s�ב>�..l�^�H���nj�$$Q�GT(��,���Q���'�޽[}.��B���r@y�MP�������֡q)�Ck��ԋ߿>�x�s�/�@^������;|����Z�e�~���%���f���tk��i.�z�#�y��g�ܿ��{N�e��*�Y2p$�Q'uom?�lè�h9��l�yDV�v��?-P�W0�o�y�=�g�k�YY��a\�Ω�{T'a��k۷�f��k��������p;�����;��;��7B0�C?ڣy�f^�"\@6P%���<s�)��h�Jp0Ć-��ؙK�l|JI1�[q�QW�x;z����>����a0R���-�~G:��gci�©]h�������� �X82uX���%tt��ϥ�o��7�6�g+nR	0�N��MV���NM�rr�f���2uH���~��w|�4���,h}_l���q��qZU����Cp��U����:~'���yOu��'�qq����y���BxJ�J�
?�XwB�?���]O*֏���ww�"|��3�V$��c��a�Jk1�A�����E������9�G]�]GǇ�jh�g�������$G_~1.�~��y�~�R&SD��m����ƀS's�6�jZ#�a��^�"7�h���a�P=�D�ӛ��??D�϶+�SL�{���d�F��<�o�ڱT��ToI��@3u
sͫ+�N䮑�f��,�Mcޝ��u��C�|��\Q���D����x���� b�f:�RO摢���3/�����ǎ���� Y5uO�Cި�g���c�����j����WUz�ȿ���|�����=z�(� �=[n��i�{�9x���߆\k��-H���r&�*S�ۏ&YL�<Q ��g�@2��`n@��:��fk[�:�xo�[�� �2�@D	�v��DY5�3 � �[b���h\4⏿"�H�Oh�
��V�S��(��σ@u.�8R�E6W�#��lE���Z�<�ԕ6^L�&��[9�zPS]���ƺ�\��)�ᑾ�7�߿ �{>���s��(!5�BjiϠ8�iVAABq��"x.9����n�a�[^î�Ы���\����N�����_"�O�C��$�F����%�myNz�70���J�a���������m<`�'KꖜL�{���r'�fwq�K��=�SIA
�~�5��u%>~4�7;ED�=#qhA�l�G���2Vf�����yP�ŉT~�ٛ��ba�"/¸|~�x�27���������i*)�6ݻpx�_Dd��ߎ;�WZS�H�LEI
 �@u_������*��2z�J��������	zu������Y&��C����L����E,�^��Ϧc���h/t6kd��ODD�r���(�f.�?~֠iĐSM��Q���hypȽ���,i%V��-���E��B�O������?z��J42.���j���i�x��@]>��h[^�r�����Z�q�1���18��0�ԮZfA&��Q���1)eX���*��G��d�UWjN��1'�yv�RW�ć`q���iI�CK�m�|+�X���
4 !vf8-�����m$j��)�f��-Ⱦ>T��}���Q)��[B8_J��4�qy��{�[6@�p8�l�{}���@�uzZZ[cVۚ'��%��֘��̿�����k����CH8ۋ��Z����73o� ]���6��Hj)����Xeq����~N���q�K�<��QFbAE�{�����M.��O>���W���혤����9�A�-x���A�O��$�#X��=�V��;zs8����h������g_�:�)��J��E�yU��<+��e���"_3ss)WJh�M�"����y�!3�%��aSo�
�.�`�{}ccg�T�*]��ڄ%�#;੟H�bG���nK���:1�|�o�3�*�Y�#�|�	���j*�55Qj��徛�A3�2v�Z�q���J�<$�,��Z��ӳĜ�$�:�K��ۇ�Kfeo��W�Pu��1��7K\���d�9��߹���ڗM����������J�:��O���N\�d|����Yk����UP�z^!�F�lsII�L�97�N���֏Q�u�.2&;��ɒ���}�N�8yc!�\��O]���%d��q8{ߏ��K0� ��Ͷ6��&�>�����W76�_�/vw+|�x�Μ��A�DW_�H�ΨN!iG�z�9
51����Qg.LZ���������˱tM�G��J�[8~j��N�*S�}�<��≵�!�؆�*F��u���x��	D�2�B#�������^2��]���h����?7ܤ�-I�8/�{D<�4�������^��F��%p��x͈{;����[|��	?M��T�����v+��������=����P�L���oxXl}*�E-·��Ts7��0(�)?y���t��rr~�c���&��3�]\�i�aw�}*/O���7N&��_�� ��X��jl��3U������d�v�a�g��������c��rܷ���%��h����bB�I}�>�0y��r��!s�/��WnG>G����|��x�G�?y�h��Z�}uHH/���������~7��{�M���kb+ѻD�ND�-D����G��-�[�&�FD�D�[��}�s�8�e<c<�^�Zs^�k��ֺM��$W�PM[���������[g4 ������kt�6�9�����cOψ�h�h�\��@'�)tR�X�if�7X2,N�+p�c��� Y^C��Wޓ��i�^)H�[Ě��	x���ѡ��(9��(�7�74pm�\���n�R�$�~������Iz�|���_�����X:
!qJ�J��,֏��2V����Pm̘k۸!f�Y���̾��!��I�L W�Ұ�S��b��I�Ќ���dM��{�:=������`�k�X�Ew,';�Qx��
��@��W�KH`��D#�d;��#L��C�Q��s;�󬽋��gZ�z�3n�8�3I�;�1;�mW>?��R�^��$�"i��pK���t��QSW����J�����q"�6+*<Z'l��`e���0���q���\��ҙ�T���G&�(ǒ[RUђ(�Ճ&ߔX��U�� -��iN�\ނ���S��b�੼`��SD�c�*"G��R�c�T�h�ݦד�ԒI&~����nlz�y���G�t���h�xң���*ݘǔb���tGg]�������#����o�v��7ˡsT�e�sM+ӌ�����ҧa��{w�'�N�bï�I6���i1��c���/�F��N~=���Kx8�?A�T �����l�������ߗ�`�+�~����;���[y�+���g��"ECz2��/��������)1�SY䐺�o~��O�}��פ�xd�z�������=̽9~����A����:��ݝ���L.o�9i�O�vk�u.�8�xB��1�R��8@���ˌ[M�J?W%:�6@7�MM��*/��:�5�7�-Gj��9({s;�'����݄;֙������M��4�i�i+�hiU���-���X�'IQ3j�HQ�i�c���:�[c/���7� Ij�c���L+0�ؐ.�0v��T3��]x������s�Qӓ����^+�Sh��s6gf�Dn�N���,�]xe�Dal<�rtûYLra�� ���K�}��`x��<�����gP��F�jλ�m�{��AKX���P�{Ѧ�
��GV0i.m���Ğm4��6��f5 s��Zl���][�O����8����ո����� 
7�;:�:��s�tv�y��of��uv�*�Sz7.�#�:C�,�u.�<oSsQE��� ����LK6GD,K�ᐓ��:�;��R6g����\����5�z�.�/�~^9mv}ƙ��ӥ�T�@����t���Cf�A�â�����6*[���mEYs󏉷oΆ����}�l6���K��5�]k�O]b�?{����oZ�q�2p�	������T��h���'�j�v^�O��2xJd���@����47�U<~2i~�C���F�lU��J��Q{�VI�u~�FSk��t�t�uG�=)�����d��X�O3H:�݄�/Da�
���� R�D5��8Gt�H�Я���\9����-��L�L����;��}!��  sQ�oJ��=up���%��2�����w� ���T�؊ê�v;��9��~��������2���=����h�`���)Ѐ��k�vt\|<Q9ɫ�;/X�xn��xkr7�G��w�I3yJ�N	K�n�
N(L��q4OM���Sl���Č��[D��� �CN�!~fi��֚4ɞ����A�AΛ�Ɗ2���c��K<�
�XJ("��v�g�t�i�f�7c4y��$U�{�/fc�S��#T�W� �g�=֋m�10pG2��_ں���NM�$���%���D�n�w4�8������QJ��ȵ�c���B��|4PȷX�|�& ԡ� #���3�9u�����?Db��_��~&� �r���I*Y�ʊ��9W#���E��n���S�Rn'��N�k�f�����P��v������$_�W�D/���0�8[�x���c5�59�Td��Ԇ��anT�v����?���ha��s�zn,z��D��x��S(ӋFP����jUlf�|�###�����>Ûvu���y�v��ؚi�-�h*?���*fi>7�V��m8����a���;�[�%bP�Ҹ��W__�R �8���p����$�}#������*�4UD�L��`Y� �B�s��M�"����[�q�KȰ��As��bX��N�EG����K�Y(p?�����۲�ɂR)�, ;"���T|D�]�?Bp�V��U�EI	7�����?�@������/��ݓ��񕑕%̶x��񫑒vY))�� m���yx�vɓ��z��쑹�t���M )�]���/fFFK��R��I�����F|��E���~s�aċP�b��~EZjꗓ��
�����=���]�)g�o�ɉ	n	F/|�r� z���o+[gm���1M�cR�׼���w�&����F�}c��!���{��+,b���e��hN�ui�B!G����F�Cz�<�C�J@��D�2��>(����h����$'�Dm@�paa�=Y�Jc�	r�O	―~����1p��C��b0KVỈw��y^��������m�[�����Q�S�o��_]�Q`5�I��r6�:�ƗL���M��3�CJ�W$������?�r��1�G�<%��lu�q榕������sˮ&!��s� ���h ��ö�N0)_�$e}5h�G��dN���X;n>.p���]����41���׵��CJ�vE���///O���q�& ��Z4�a�n0����~�@@�����G;�=]�;�>i�B� �s�������N��_NL�Ȱ��P|�*G�o���*-�x'CF^&�-������f�b����/�bwd�wvh�<2��-��rۿ�Zߊ83H0���<�9�`��0���І�~=��wvt�֗N�s�$��Ls;l1�7|������#�T{X��5�ʓ��i6�D�H���5	�M��ޅ�����`��KX�jq�u@�+���P�O6$%(i:��n	8|����ǜ+f�v�u׆�䤘����nm�n���z�#���~����
��+n����䎊�''��ι�{y�F���9�&�]X�v�W
�0 ?b�(�
���`A�W#Uo3*�ڪ:�DSK4�J{&�sx������wu���k$��ro��h��w��z���	H��:�ߗz,�� �$6��H<�>ʴ����r��!&�Ud�%���Q0�oo��آZPa���C�1�`r򉘌��-�p�q���l���ߗE~o�|�<�Ё4ޣݗRCSs�I$���o�|�3��V�XV�wK�4�j(e���u���H&��Y�n��}7퐊�.�R�#�}c�v^!:�8}����8�&�e4Ի�o�m�U��B��-T�"Uoc��(�LIM}�N�]a��[*���fff���)
p�nˑ��I*
R�s#��$LR/
K�_��,�� ����� �)�c�QC#N�"
,��"�S]s�3����Xݒ�nnx̴_�'_D-K�����ˌ��2?�6*�?k�h,$*:W���߽0`�C�mF����G�9�]�pg��A���۫������j�G�s��B��Nea��r��%��M��D>޷
t�FmH�c�ٱ�{ˌ� ���T�v���У����cct �������L[s����s�Ƅ��yU�{&�]|]
�]�����@�K8��1\�oW�`.��������lL�b�W��g�M�
��hL>c#G�r��{'�JJ��h���7u=�o�\��x�,���/XD����=�#��˳&���M7*ߥXMx�HC�"�g�T��ERcF����|���w���T���U��夘e*���R��a��C��]ϦnB�	'�y�4�_Ic���K�x�4b�/95�'w�-ڀmLΑ����&1X�j`�#>���ޜ~�ez�K}��%�B�b��ȵ��(��^�(�_�'�ݹS��������B��`T:@{	�g��Z�0R�im�C��sg
��c������` ���@����#O���m�(.(����|�nEz��*�6f�/�v�~��~���������M�Q�����KV�;+*�x20�?�&0��Iʗ=X�n�j�罯��,���Ƌ��1՘R)�ć��>��ݳR"溔��(���R�O4>��2�Kd��~c��a#�fUX͊�?'�ޡ9܁daN��r2a��4���C�� �{ﮩ}.���v�9~G���?�;"�+-�S�C�Qp��,��C����o��k(2��ܸ��}�]x������cMr�?��l�G�?VZl0��ueD]S��\��e�փ�P���W�O;/5Wd#����7..��IH��eE����>�ԕ��nN7��+x>�|�{|o����h�ܵ���w�ܡֳtY٧k��s8;{�W��H��԰"�r�{��+1�B<D"Fi�?�*�:z{���m�}�-|0բ��ՑZW�\�%�m\&�ø
D*�4��kN����G��i�=�f-�:5�$ҳS�S���y/�B�9���c) |�bꂕw��/߿���8�:
��XQ�\V��MHȓ{`�������S�����ݫ����C+)���&t���u/���M�UKo�Ͽ�����(��~l�ٮz7�n�����ѳ�f;&{�+Ū���9�(�okk�5�1���VEߋ�^���z7�Y�8[���3��140j�G4d	P��^��w��XG������S5�����EҨ�1�$_cF�d����?Ժ6���{�Ux7|å��^�5`����X����[�ty�4��݄���_Ye����J�.?���,z��h m%����%1qq2�t;��¢9�]��55���"��b�?~�4�6$�b�^�����rQ�~_~#3)A?�r�Vf��2	/t�֗���M�놡�YX�4z�X��RT�	HcTrXD�o����p>�t'zIN�wǗ����`�PlZ��@)$�3ٹw� *���O�	�nl����������\m��^����rj}dXD���Ѷ �x{pfs�$�[$i���ݱm��O�Ē��ɔ�����Q�m���'�,��Ճ�����x	ʣ�?JP�y�|wЀ��yڽ5({��q0(��r�ǀ��H�hH�PkC��1�=+���ߋ����[8[ϱ�ttH��#E)�0�G|��= �,W���y����=���}���~Q������*�r�֒$��Zq8�Q�H�\L��e�l���8�"$�5�ހ�������f"�����:�o�1',�I|������n���O�%�_+�3�Q����;G�������
!A��d�>��74"O=<���y���ku�'p%�/{JDQ�_NS��8�7_��h�=1y�@�q�w�Z�� �Y>�g�s9��%`�Y���<mYW��P�/Y����T���ҽT�5��
��~�G	A��8��߅_=�4q���]�ϧor���i0�[LU)x1�{��S33���jf��^�6��مȈ�uG���C�/+#K�z5�Տ��K��v�Q����-���������vՕ�R���GU`��ݗ����>�vc1Ak�)o�'�58�I��ͤt]�c{܇��!��4�.H%r'���G�@2����[��o�����۳��
��Y�Y�$��kbt��R��{q� $SU���m���mւ�rr�o�%%p�o���^Xu��4�����z!��[��-��-:%��2���:��=�+�{�h_���B�3��%m� "66�~�\=3���s$�Cb�O7��l�SA�~�׳[����oI�Q�JF?^�Y�����"�6M�\���L��省���y����j��j�d)! ���O}��j�沆������cuEʉ���"�5��|�[�Tnk i?���k��^��o�ς���[&�vg[q��Hh��#�k���MiR4#C�i�-2�EW���	��@w�<�J�h����\%��s�$L[����[y�BO4���u�ws���3���U���@j=�����S�Q�/�223#���&z�y���XH1/I)(�q�»B���#��������ZL+�C�|�)4`f���')�R'���XG>�ծ'p8X��֎|���_z�M�H��}� ��뇕�=�i�T�Y�8V=%�(��g��ZEt�C����ͤa�:�S�G`a\V���pK1/4/O>��8u�W�;ZW�{Pt6�F��}0~7�¦mgxuF��k����+���I�8�NNq��Oc�����eC����n�z��?{��x �\%��z�
�J��ٔ�	�]�*�����`�i�,�dƧ���ؒ��f�ݮ��b���|�#�"�B�1�0���S|D��:Q+&�p�K��J�v�}����Nʫ���/�6�.��pz�ϝL V���{��cw�fׯm�۲ӼO�W�qk�uqm�C#�휭����P����`��-鬟�������+<��8
�����JJf�-U�0���<Pd �&F�}��mr�����D	�~��f8n9������1�V'�n�W�i��UZ�!6��K<s �d(v󎌈�>��YX���u7�P��^6�@�^�>$�B��b�H \�����CCP�!u��E��,�kk��YV;�|�:(TT�	�:��íYaM���'zt�--����q�zh��SB��'�ij�U�?;�׷�+�
��Dh �xJ�-����	r�4��+I�3*�A5|��!��5aDR�H�����~r K2������9����Y���k���XŐӁF �f9|�č��Rvl�e�0/hB�����ID����a�ũ���	Z���S��Sx�V�-62���2�� '�=�4y؏��H�T��_�3�p.�B����4t�z�V���.3��O�]�����Z�I�Ν�¦�4�w��D�B�w$4��'(��j�"�5=�K7�^��$��9���ǾvW�w��ty��E�(U��JGĬx7;1�B����5K��؁����G�`�g��@.�ly"�yJCc�\�yfFoa���|�nD��/�.�F.GQ�&+~�P�:�X��|���j�Wpp���Ы.2$\{1��(9L/U��3.����W��O�+X#��B�*D��S������x&�ge-��n�<5��ǋ�>Zƴ4��Y��L��0��i3�)P���5D�^B��@Ϣ=�Gf�l,�|�.�VbB"*��^�vͅ]~S��?���2��@�f�оѿ{$�e�߇�BC?��k�|�y��[������^�4����Z�0�W�&-Q~_K�U�K���Gcﯛ��M� ��D�4��qr�7�\�^��O���@(��H��쬼D��}�+�$�srq���h)Ҝ�;S�^�,r*�8ON�Ґ���"���{�ѵ�7߬�A%��-#�������\{k����Ɋa� ��`�3ӌ��8��~ro[Ú���bZݣ�����6�>�FYޝ�>�RT{j����Wȁ��!�'� r?��v%�$r���L��F��*�m�z!Q�����7���������(�)��V#.J+oo��B���ӧ#�Q��W�%�ۺ�?�>�����ke�F\||�_���֐�ŚlAK���Hd�Z!oi,"kPX�k�O�������F�
��n�@b���=���J�SĪ�ȭ�����D8���g��(F
9��[�v0}�&�����mё����G?��*Ddk4��(e���3�Hd�f�w�9<�m�PX� U>�;a��Y��ΐL�@6z�H/A���$��K��B�Y/'��W�b�=��R��mR���M����V��Q�ּ�?����0��;��ڧ���~�7�aig�d\_�OC��W��ŗ����n	��Gc���X�����(5~�D�b~&X$65��FWN;�阱|j������QP��f��vr6�/�{�Y e�2g�}Nh���c��G1������z��m���u��4��«��e��z;7N|~������ U�mF��4���Q読��j�A���3J~��t�u� ����(���o/":��#N���
E�T	dNxP����WRP�GO_���MW���{m��X
p��U�O���tq���ɡ}�7�/X�J1A�#�������s�ef��I7�F�u�&þ�c2�sw��������:5���:���O>�(%���Cc�SdF�������Y�D���1ǺR@}#�����JJ����@���d���[M�^(�Sfo?��ini��O�͝\D@EPh;��]��[�_J�Y���\��'O҆��N��q�a���D������u�ua�K�� #�Ao��| ����l�	x�]�W䙶02����Ä�z�-i�F>%6��"�y>r�3�v���(;t��?k~|#�V�5��H��L��8u\_6pR�^9ZU��	؛�,�J��sQ��� [���>Lѩ�&,6����&ѵ�����u�ۦI��l�P}�	Ѱ�M����*eY�nxߪ4�kV�ٚ	B�	 ez���@%��$:����D7��t�nnH+�܈:u�5?j�ĸb���N� �ؓ�?h&!Ē+�7e���B�ofvU�!)� ���f�'q��v�y����PoZ����E��޷� ������ö`�Rt.�q��a����?��8�����|t��|g�g�f^���3Ms�$H�<����D	Q~�=ܼ�C���
m֍�y�e��4��@�)��=��-),�ظ���b�@�B:�cR��w��G!#+��������4O;IX�u2h�_��%�ܖr����=��OMJ��7�y�ɋ�J���Ò��v��6����4ޞ�FA�<s�*;þ/����>���k�R@��p2����'wN�lLC��])Z�`�F4�?wd�^�90� u����m��>�#{�4E#k����&��֗����ﰰ �_�pU)��77#֦�E3e���ð���ŉ	r4�_�z	Ҵ����pd�M��5o����M@��ܱ��(ƨ��H�_T䢬���~�/�/�Ș�2ܔ]k�9���J��-kW���Û�T��rE��>o��J�q��� ���L�UkAj�xziY��I�q�q��vG#��lm��%hy��s5�d�}ҭ����o l����%&Z��0�E���xfvV��*lA�#��Q��`:�	y�e�h��U>�����V mTP�$w�E��-�rj@�Z�(�O�;�Id���֯8d*�ӱ�[TK�waU�_|C��G�]�����1�0)F�J�;��&�c��]�ȑ}��Mr��J2*��d��c����h��"�,2fc\�P���'��<����#����R���&+\��桻dm��kS)�J�����O�s��@��JV�o��>�D/8�������ml���{s����^�p��eD��9�W�u?u��f�tÛ�<�?p�<��y�81����*7�k���rȠ���x���f�3���]�kH���,�r��XJt	��	����������A�e���ɴ�B���Psv!�N�	�DOg=��g�̏�����䒃T�J�f��������x��g��U]��E(��o0�D<q���GF(�F"���2||�Q�r�O� J�D�g���$%{�j9��0�l�c�\Ůէ	`Aً�O9a�YK�.�*7!�KD#�����&��e�3h�إ��r".̾[��EQaa7�w����	6
��K[�At��e�����i�=?Xɚt��᝚�W���ec��ϣ������A/��HJJ�Tļ�޸��"d��=��߁;PO?�I��P��,js-��I��AX�Է�s�.��KJ����oƿ��wz����	��%i̾�� C_��hr%(�w��/��4�EE��@A��&�:𷸟����P�k_�t�2�I6�&�۲#���9$+{6!#�;W�󕡭�<T�'X�hX����H5	�$�dL�}�8�F�����q�k�|�:��S��j�h�_hQ�gӻ���@��~${t��������\ah+�`�U�������;��5O	1�q����k�?�D~i�V�}_|K���߇e�|i���XevKmaG�܆�vב���<��GG�}}�I�R6&i���ڶ���:�y`����@�A�@g)2��lo��2W��qUm�X�o2�b�h��.ہ�R��>G���
���#�~��}R$K6�am@sc>�*Ж�OM��7��(�I&7T����X]-=2�	KQ���쥆n�GZ�q$v��$4�1ęu��R^��G�c ���sB3�{Cպ�n1	�X��N�}�%��L.�q>��b����N0�����lY��ɨ����e�^G|����c��E�n_(��aUb_�"�R=	����fc�O�f��34�FmHc[]ň���QKMyz:>.9�=���8�>|Q�P�7��U{�-}gb�{��nM[񊹻�K|{<Y���#�����oT�q�MO3�S؂�J��$`�����]19>R�c��`�L}����,�`�'�/�#+��G����^4>mfDf�5�.g���Œ"h]E�l�OE����f�5aqP$,�j �6úc����S�Y:6)������<I�o�;9:����4�!�WC8�f���?/i�ˤwG�Y��Tq�/`0�s�=_)߳����i煱2��oi�s�@���G<e�	|Y����}�r��`��MWW���z	�ck^n*+SSR�|�
T���Ǎ'/4x��^����O�t~�|V�q���ɞ�q+9�*�a����Gl�������!��=�fW����@�c)y9n�N�u/�0@� �G7�|��m������QǺ�k�Ƽ���B)� ���Lѫ��Xc_�g�0��fY��|)�&��w���3;v�p�*�p�^m!�,��J�]o:�����Xw�l/�Ј��� �y�>�N�ƕuk�%�S8MAs��{�Yf�WNBП��������KSb��^���M��MO�Ɂ��ŝ}�?�����H5G���$+:ÿ��P6���Dr�2z��ѐBw0���A(a�\ ��V��c]*���/��:	�b:%��t$�s�x둝����\�;�U��G���߁��y�������!�'7�\��fh#Q[��ve��j�!ܦc�h�ʲG��D��	�����)]I»\��������`��ә��nړY߾ 0�96i����I�R���tE ҥ�� 4T�a[�+XR� �(IѲ��㣵����8����"�e��C-��5���e3l�k�Muj4�����cy97tcek�I4O.3ytOէO�w(	�$$>]y��91IIa������P��tшA�c##jNb�+c	�ˀV]���|��^�S"�� y�`=S�z�w�_�٩��</u�B�)�K�2K=��'n0���:�:��.8��"�΃���f:�j@n���?P�L��H�����C[[�w�<24��'�D��2��xY׮&�xD"ɝ�%�;67~A�̠%�=��y�8���I��Iu764tLֻ�B}��Ы�A3���@�,��pȊ��Y��DƣǏ�
Y��m��댾_��Yɦ��r�^g!��T����265�Ao[���4�iD.�t�O�(P������C�RN��#�~�Z����4�$�P�o�V"���m�"`rg÷bw��1��!�-u:Z͵��#�/#1��{f������I/0���5�qm|u�K&��_�� ���?�E�����A�.�Zk��ң�#�`�)�YC�6����5�>4����x����,66��"�B*�Ĥ��+"��Oq����t����t�%���7� "	a�MEZ���!���T�5)$���=��10��z���Nߥ�����tm�֪����p�Yォ(_����^v�ڄh��ީ�:�EІw���pQ�������*>�|�߶ߍ��FT���5X<���H�`���J�k����?:~ed<��Y�%��?0�3ߤ��rlL�0�yt���������] �?j�|[�w&6I�,Щ�g�O�dH���0�)O�)>��0�����g��8p5DRC������3�:x�h�/p����aqnBC?� �ߊ�/z��~ YJ��J�����:��u�#"���<�.K�(��cZMI�Lc�ZN\[AT嵭����
,C��<=��c�{��xn&9o.7u�2BY���\4�����?_`#�ɑH�cBa�^QwZ��3[r?:_��*�1�<��f�7g�}�k`YRn�����{lB�1�m�.�w�L��l�h��9�V�@���
[�a����lƸ�����G؛��楒�]\2���4�4H���-%��_�񃢑���"riO�bJ}޻9��S`�<�ώӞyy�$����A	�i��=%v�v(�S����]f�ꊡ�2�޳gϢX%���t����*�\\����p5-X���s���^`P�,}T��fZ�)�x��������qz�x�5pS��|��1��������� %C�	: ^�v9������=��l2��--�2����칛�y����C��Q~\}���ǚ�9<����t���������q����h�>������1|��
���^� *x�T���D+�M��^ sO����������(���j��k��{JM��@] �d������ma���XX�;�;������A�]��r ,�oơ�(��T�?��`7�+6������1A'Z	�M�G&��2!��{û�K�^M��u�v7%�+�gk�����]�ul�z=��Mz�R�v�<Ffzu5�w���>̴�N[��D*�c}=����%yk *gs
��\_w�^#�����Au�io7fNN��K2Y$��"���PM��k� נK���N�+�	�-��M>dުC�tDP&��餫�¨=B��ˣD�Ք��'���>��ݓP��P�]�]��Cm��kfC$Wm��c���(�q�z�o"�ڍ�<������l��Au� �aSkJ�Xaaủ�cyc+#ǁ�;[�e��h0Y:���Ι��d�7����"ꊇ��)�[�R<��3��ܙ��\�:����o�r6�A���n�����}�t<��'���
�hܮ��������g+P��x�5/ҚL����,�s��cwH7/�Ytd��0T`oH�b�|^�4O�\�N%�J��<���G{�\Z�6sMU��6n+����N"VPK�l{v���ɶN*�_1^.��(+J&)�kɪ����;�������n�qA9�p��]E�Ũ����⏬��}4�R����wa!!����5��@�h��E��z�A�E�3wnj4���L�Q�b�?��ገP#��D�g���w?v���y+BR������uT���Ń�X%_,��������3�v��?����h�N���Ŷ��1���p7/���NP�B���5�#�WQN��D��ߜ���2�B��y-�����'zT&h{ěۤ�r�N�-k4����y�[� � 1~�/�7ʾPc㪴}��"H��R��A^Us��.G"�^ ��=�:#�	��uV�Þ�2�T~�t��簳,�0�d��uLE�F�F�[���wI�(�(�����r��� �F�u��he:k��8�O25/!KN3�{�n���>2K�g���|ӿS-������1�^��6wת^�M��>�O�^k��,=��i��Ͼ��}?�H�@�~����GxW�����2�hr#{�1�)���^I�<Ylm���fXN!&��"�����Τx�=u�%.�9�k�Q����Qd���C���F�r�����Ų��>Ǌ�[�e2�����D��]s�,I��W~��Hw��7�����)$@�0�)�TF�����[
!�}���F�N	���R����tO���waŶ��"I�:Pu6�w���p���>��l8+��M�*�+=+9�i~-����;��Bf^2�a�%������V���iNS�9�i��ޞ����Z�x�"�IKQ�e��M�͆���1�ԮEnb�yЩU3x����HZ�ظ�,�n�d�FE��E�v�V��IC��T ����l���O}��7���Z�N�x��W��8�k{v!�<_8����wP)�C;��BT�P�Z-���ocǵ�ܓ3NJ�=��7�p��D��V~�,	���w,Z�����{0/�O낱|��������<{6G��	&��(f�������6�C�ze��H�%�FR"< ������A[��b���U��7���j�y�����ꌨ���n�z�!E;~�/)�e�������|��y���,��ȭ��$~k��w���h������zM�H�^�H\yH�gU�UX8J�i�:�lH�do�r����/�F�.��s�_�wͿ��7��:�v�c��i�4�O�#��~�?���](%~:���#t�w��;��]܄�K���#/�4.ѿ��Fq#U�[W8�����5Qq�}��M/'�1t�l����g�wN�#����vv�3�"Vӓ���/+F7㙤�I��x�����K�[9�����,>B������3�3m��f��;����W��:{� OV��k�z�O��Z�j���� 0QK�I�#�+&��όX2����70x��YnҸ�J0Yz���қ�a4�C[�.�;*��'�A"de8(2 �($�nOk h�'���t�P:�����₠/FO�M��s���)��6����eNsN���H�+����t �Un�{���4��[�u�o � <�����Կr�/ٰ"%#��ޏk�`Mo��ӀO�Bwq�,�����"�s�-ػ��赜�MA�J&�d	I`8�X��ӗ�1��5�p6}�0t�`�ÎO�7R�#}�(����K�(Ⱦ��
ߴut$���'�,�FWXD���e{��}�v ��ᆔ�L�@�����B\l\�����֡����q}}}u��hccc�'����˽}}Y<I�s;��p*���8��,�%R�D-�;� ��i>�5��@��Nwx:��J��772�����B�xS[�����$�3��_H�t�&p�y?��Rґ��qo��~m4�y��#}̨@�S��PB�]dn�q6���)��� ���x�iF���<#�C���2�_��W�'���2�����W�t�ᓌ��LNN��>���b��[��YjF��-�V���զ��t��k��i�s�*�6�r���Śbz@oN��
8�T@k&��d�j��XN8GwB.�>-���umb
;
�,�:bSJ}�֡=�;�+��0�Ww�T%�*ec���}�!���Df���[���/�3R��9���W�vu�:����ۋ@�N#Z�fڂ�4<�q֔����|��*�QP`5	���Ҿl&H�ΐѕ�J��Z��'x��]'��(0��Ug)�A�=�n%����D_!+������0-U���N�E��,̥��L{s�?�9����tm89e�Z��5!%�,!�<�dl��b�X������u��^ǳV��w����X��c�'j5X쫙�����?^;C��䣷�W�x�o-����(_JA�f�����a�`Rؘ����ޖa�־�!�X��:�`���R�*�jEB��5�I�6"��n�x���7g�,CB��&��*��X��##���+82��MI����`F�'���nQK�,G�z8q���D��7t�-�v����űc���}�(�7n��R�#���o`�>imj?�����y�d��T�̵�~��y�J��g%z��^��J S�C^�9Z�~$��"��2�1w`te,��Q�Va�3�a�x�3X%��}r2iU#{��&��>$�C�cza�����ǁ��7��
jV��S�X)	�lY���;�K��
ᔕ����s���p~I��X��mk�vP��20@�������P3u�?���.nQ ��I��Hcy&��	:;"2���փX��ӧ�u���r,-��r�\��cS Y9�"����1��J��7�'7��������Ve]۶q*jB�@�|��*ҋ�r#����%h���\2���� 2Z�ɵDi׿@'��Q��¹�lYkW]3�c�����'w�Ѩ5/�Ҿ���G>U��;�J<�^��RcKӗM&��Д�Ԃv��>�/kJ��eΤD{M9�&�~,/!�T����/��`4q�p]��R��o��J���gn:�:D�(�=����C���&Ly�Id�����^��O��$�f�hL��}k��=W�,)\�	lT �db�%Qw�{\�|�=�s"�4����Q=?z3��Dz ��GC�6���K9k�6d���wH�c>��$ߒ>s@�OMA	�^�h䫮&#Ŗ�����~/i5
������W8G���pI5�����<E�i-"ݶ6Ҡ��E�wˮDV�Û�ßX�p?��K�4���]�5��-F~�mF��G#5<�ڂ��b�#)���-s� ��Y���o:���5�J��iSG�b	��D�u�Hd�`�#c�bz��޴*����Y掩)�E�:��A�pF	O����L���==�P�!�����$@R�L���TdUӟ��L�f�H�ݞ�ꩍt�^��(C�p�;�W�`
�Q ��3�C�U@���[��tK��'�n���&j��sGDH�ކ]�v����p��N�$�;�Ǚ�\_7��N��&40�S�R�Ew��-�`�^8�|�~�Att�H�����r���ǖ�-��-5����iz�e7����JY�r0=?{�#	�EU|�=����H��wz�MC�m�a����!��v��3ц'�v�M$�R#�<I��M�	߬>^v+wqt���������/�|��XX�.JS�e���@ݱ ����hAV̻T�P�l��.q:,|TY�����ܕE�N����)R���{�=��5�W%�n?�)QZ�����}��m�'�NQVv����ݦ�蕍XE��\	���<��k;m��4� ��]YbɄ�盽B��l1a���J�R�E����dx�[�i���%B��V�)��G���ל�.�g~�e9�xIH_��}��d�__�"v�Fu�#�X8��q��w\LU�����G��1Ҙd�\��F_@p%Y��x���k(��Qy�8kr��	�)��7S[݉7�]aʟ$2���P�5���Pu��T���?""�ұ�U�8٣8�3#9��(�H������22BV6�J��3�w����?~�[�ԍӹ���|<��u]�Wγ�ַ�<ob'�vF+� �m�<�k���R��@ʝ�:����"\Cګs�7r�X���*C.6�fN�� y��l}�:�IO�S�2o����R��F!��ռ��Q@F⊐�u9#��F���hV�h.�K
0Y����V�)�V5�_����%��O��3t͏t��q<ڪY=��c�#��-��gX1���V��w��P��2�����+Ȼ�z�	�>벢��z�����[��I�3��{@{څF��\�(�I���y����VYuh�����8��l����J�Zg+^��_X�1��_= �
2~�D��b�A|�̢�[�յv�$)�ӬXOㆉx<w��e��)�4+��e������W���uiV���[&u���Ra�=,{(���'jl�Qe���kn� �������%ý�%�t�ЙtޘC�ﰹ�z�,#ic�73�u*��e�-Йtv�!ǝ�q]8I��L�F��v�ߑ��y��C�E�����6�P����4�Y��W����)",��L��t�Y?��[!�$����y�s�8��Wj�]���6�њ���RKU6zѫ.e�)}�M���ڕs��X��/�;}� V������m�߿�KN�=緍Cb/�fЍ�D�_I}x��K��J�i�y���tŘ�dt����)�S�*f�G�-܄���P�^+�u�o ��;��X�$������#W�-�$�����͹�\���;.���ƺV��٬����z�/����"��4*����$լ[n�X��h����Ak��F�?KV�!�q'1���P�+��*C�"��r�6�����2Z�� {�cc��s!V�OB?h�1��I/�#��}d3�/g�`3��N�-��;ԏ�N.��E��a �$k�t���R>���Y��1�2}X�W��z�&A���ѯ������tҴsmOr�fi+V�^�B"r���ik�ZHɩ]*���;#�~�GS`�swY-;mHd���L��d���n5�Z��=[[(벛y�>,,�X%]��q����[y����irE���ٽc���9��hJ¿ou��b�Ƴ�m�c�
��z.V$��~�D���Q�(�F+��y\
H�X3����{0��p�Ha�snW���h7���	G��Ɍ�0hJ!
j{��_}D���f�<��f
�V�s�E�<��u/^�3��o����:u�}�����U��ޑߏ��t-�+�=�'�ҿ������d;-����n�9:�yR�뗗��Dk�+�ѧ�+$#���D$�j�Я)7���dYu��nq����W�A�VF�-+���cP/���9;\�S%j���|���&�Y�?�X�O3a���'ߗ�I�057o����6e����}�n�JnM�� ZG�	T�/�Ɍx�F�3�4�fOڀq�(n���#�5<��$�F�k��~��+iLV�W�����V\;�)K{:;-����z� ���`��QF��u��3 ������ɝ�o�$����t���d�'hTX��nI���δ��� ���]�����GT���O7���M���5�|3����; ��<)�S��{���u�2��nթ�l	�����s��|��&��T��;����j���L����ҫ/�2���	�ͭ&R �����+#��x�e����ڢK0͊�b����T��h�K+PI��S�4�׀|�)���"�m/1�H�`��%�>�_�㭮hg�I��klW��I�ۅ`��@�S�ݢC8��N�o���m���L�?�������{!�Ҁ�z����\\:	�q��f%��ȶr���]CP�.���!�0	��&$\6�k� �7up$J�׉��Y�����'�`.�����gS��%�'��2��?�D��N�Y?���H���?;?������m/��G�)��X�ʱϏn��]�b�|)�}��~��E��v٤����c���+��F%#����i����ۮ�!�I<�h���5N\vְ�>D�P�z_���B8%�eM�;�����r2Q=6�0��}	+8x��QGl�`u���NB�͗�	>&˘��A~ͱ��Ԟ���y�X��e�]i�jo�G�[*��-π�a�������4tZ̪��R�-^�����̩y��G���M�B���ʂ�Z}aa�l�w����e�n����'��J�C���H$�TAg^�]�~��5@w���H������w�sN�/�L��"ږ��iپ��z�7����3��^i���H�2�.��aD�t��#�ҟ"��k�4}�E㕡��7PI�
5f�H�G���!�W�/��Hר`g,�������hX�=*������V�hc)�F��_�grgU-����&k�1�{�	$iؽ��3�0i/W/`���r�C�4���A���&� �0���V��3ir۬|�@����Is\o��T���3�6�$�'��rzl�X��8u|��߰��NE}�
�n���2wK�Jt@�+�3\���쯨��IL��w���N�c�O�G����G��Ľ!W����cͭ����+JFn���X�~�W\0����EQZN�20��j`#E�?h��o-�-��DSL�|�J����F,�	����;V�m!���b��}\��fp���ͺ�)�pd�ud�+�c�g/M�e�
�I�Ubo����M��}ۄ��\X(�(���X��g]��]~	����ͳ��KM�iΣ�o��Etު?g�x6��p���E��W�g+7:�;��><3���S!�t�~�p6#bFjj�M����
�Uе[�m��j�>~�حH��߱w�@�6S9}V�c��҇~P��8��e?�2_P��4�[2�y��aB��ƭ���m�D�7H�lJڹ�>}���6H�kƍ�\�X�t��оTފ��ă��6Nt��J���X��M��7I��$���E�T�+����k�%7������~Z�\\���>`�V�P� g�j}��X� ��Q9˒ ujW�y�;�W��B�*�@���`���_Ǯy��2}�h{bD '̵G{l�:Lsp�2EHo���{6Gk�]�d⓻�29�ႋ�{骏>tdg�F,d����:�wչI�z�ϋ��u
��u���uNQ#�SyB1V��!��c���8�j	Ų͍�[�2˒vrw0A�mq����{�^�ƃ��]��.7P:�`{Ȁ��/�my�|
d��߫Y�,l�-���2����!�V���'�.�L�2~���
==υ������ �L<놖�7�ێ�6�$tx����c*A8���!dݒy�)P��#��pI�RAc$�Ї	�Y������&��e�]����LT���<�C܉�R�9�ߘy���^F�'�G �#�ق\|Bm�9�:�ӟ�S7��Ҿ_`�TX�ǡ�~�gc�pE�s�
\Fi�P#�uA�$@y��W��JF`O|�~,�>�Z�����9����2c\��X�r�t�������; �UV	}���H�+�g����z-�����B��I���^1v��ؽ(�=���j&+v��9+�ܫ�[:���$��<�s>f�����?I�߁��vx��7Dk�.��7��}�uI�rל����`�nʛJŒ*_:� y��͂����`��ۼǇ�{z3���Iz�$�yX�ڀV2�sv�	:��=΄���(�M�Mm��B�R�kAb?q�ċ�����3<4#��5�!M�KI��N���.N�����H�	9A���0H�T1�=aX�����v�魼A�?�5�qwQ噤�II�W�x�P���e2�>����XA!2�yW6�/����s�d޽�BZD��*�i�H�S1�1/p�/�
��+����m��;!�V-���b�p�N��*׳���N������P��C�^���O�5��,�->�A���N�x�F�����] �|�τu��K�i��^X�:�e�Tl��,�z����"o/�y3�r�L���.%<r����r����&KM� ��n��S�M̶�ir.v��qmT[h�>�<	���QLi����i���EFYי�0m��ؒ�nJ�(�Z�*_��1 8�*	�&L�X�i[�W��бe�`�>{r���Mi��R�� �K
�*V3崜�1g1�B�{�5��1Z������Ug//��G? r�M�����yjʚܹ�0U�QT�&S�E|y�='���D���?�c��MZ�)��x���q���c�ǼL�;*�n��mn��${԰7�24�XYJ�?%�r�T��2	3�":,�����땒�E�@?��Γ��Qg'^�;V1��z���ݟx��q�T�ʐj�����|Z/��2� ����������P�"yHl2iJ�و�h�:����|�D�@����E���I0��cP�`��ڀ���]��`�q��ɒ�ڞFC�`΁�U��W����m.�ۡ���/iVv�~=i���S�F�03P�83�*�֩���,(�B񬻒�)��Kߍf
&����+z�Rf��fQ��޸���+��Z8����KV?��g˭�f��^ '��ʍ��u�jMѢUb��X�K"������l��:2Q-�StYBNꚺ���A���
J������bx(�����嵲B���9��馐�]�=�^���W���� ��X�%ɒ�U1���.�/�x��!��N��`���Y��E��|�_�Ы�Y���G ���+'A��ȳ+,�*Q{����a{J�ǚ�ux����a��vv+#
���?*q0x>F�i8Z�N=�\���r��`���E�k�+2����%Lt��W�̈́g]��L����.�?Ҋ�4��s�[����hl����[T �O�����1���w�����a�`�����Z��	��\� y���T�g��G~S��ض������/����6(V��w���.�E}�g#��n2�4� Ӆ\�5T�j���;�J�Uk��;9=�J��O%[����_�#d�6��[<'G�j�L����4��+P���z.�`y��"r�9�ED�j�Ɂ�f��Zӷ���=�����0���_\���M��|]�r��2� n�B-]z�U����������#�%�xr�ܘ��whd�OJW]Fy�}&�j�g���R����0{���Ot���9��2���6j�v�_�y��Eͫ��\0�s,�暦�8㳄<؞�]��^`M�2�{����6y��e�nH�]�������ݵ�w�yi�6w�F�@찕]���/w�����,b]��GG��'
�
�yՌFkv�~@� _��>�*���O�ʝьqެ�����^=��`��Wߚ*�v��w;L�l��.�2OA	�9��͈xl�#cc�I�۱�x��>"�<����9G��Vo��O���a5���ӃĴz"��u�ܕ��mDG�k��Q����30YJ����/�}q�5O�x�U�S�R�u�����.H��ѿP�Ԍ��hu�4쯞e��0�Pף�����L���q��h�M�޾4읏lȝ;u�ե��Ti���K�����۔�+?]��!}v�S�rNIXe}�eS{�_�������nwF���<��͋�������e���P�{i�D�{�e_�P�����c=q��;A��9p����z/A2�\����rz�Pc��mRc�|r�ax�Y�"l��w}��Ŧ�m����s��8���v.%�O�F�.��'���E�d���2�v�������K�rZ .�Z&}h9Mw&�������!颹 R
Z�¤�М��Z��(^ �C�/
�g�N���-���f�]Ÿ�uv�=��ec�������˿����Ț%kP��W/���юsT��n�ۀ���fP�����n��J�H�q�u��G~h$��:r� s�����~����3$�Łb-����A�����̿	���׈*w���M��װs;mZo�%j�Y�ԑ�:V�	��J
D�dO?-Y�����jiC"�3cw�|�6��O�/,CY�-X����?����h�������"Ra�����
��"m�%�^��߼q3Yږ�g_	���-�ue�^�TW��dӔ��������8&Id�bA��_�U·����h̃7��H�����=�2�����ꠡ#�uoh2�O��e��0�q	5N��՛آbڬ���9@�h*��}�(*�����O�g=��I)��&M��p��FZ㕉!,c� �X�q�(<��D�~�������nE�t!��fǭ�y�1��q/�,����]?~��bۘ'̿N�]�.����ej�r˰��|	EG�x�؅,=�M�,���\��){&�K��[�;I|.�4�W�H���I	��MM�q"
�8cv92��A�ߒ�v���|5{�'�o�ԩ��x�$��%%v�����!��g`66>�~ν��´�e�b��6�-)��X�1�)![�o���y�=$Ĩ��?���J�d���u^0�����7��)��9ɺ� 8��:/�
WW��r��p�{�MQ�����h�dL�t>�'�����
<P�}��$�ߤ[$�xՂ�E�M��� ��Y���I�.�-3K���Ei�`�-Dy<��RBvnmw�M��E�&���m�(c�z<�w]Uno������>�.뛢M�J�H�v��,��.K8��h컸8P��P1jRV��+��^Mc�˲'A�f2v'�sN��$Ф�?D!>�&�o)ǯ�脗�s\�a�������ܛ���(�|�~&�~�sl-f�=}~J��'������4�4��"��o�=���*�ƨ3��>)�*�f3�汌g��G"���`_i�t�[)��Ő2`�O	���e�A�������A�������Cƅ��s,*IW�x�,��YX���Z�e�새�s�2����@��VAW�e�b[U�A�%gkiI�>��7��:}���^Ún$�*�Ә��7~Pajj�<wh9�o��ɹ�����Qby<Ww}`��0/ҷC�z�;M����(9)�����W4+nXB�쫦ᳫ���#�+��.���➝&�y�A��'�k*������zپ�v{?�����U����jS��ݽ�/�W��7.�Lr�1�����w�G��e����_-
X$fda/�d6g�ͮ`������oy*��hp�u�v�;��n�L�%ʾL��zy��q	>�:�~O�����9�
g��/���a-o�������nb�2����su��"�`!uַ�'Iy2>6�-{"��P����^�N9<wLjh4�M��s�U�"�_��V:G*au�� �*�D\P<O�0cՌ�x_�dо⧭(U�b�w~[�s
���X%�z �齱��H���H�_ׅñ��M!t�yt�ꎽ4�3Bgw�eJ�I+E��,8�p!{�l{�{:���d����@�Nq�s��GG�����u��~�C�=�m�˲�!���L�ǐ>�;��B�NK��ٗ4]c�-$]��א5��,&���ˈ�O�����ޖ�}A[_����%�WW��1c�|��`��W��&T��[ҽ߻=�����}�J')s�<E������K�-�Ejj嚼�Jc�lw�J�߿�����u����&^����5���g�0w�GS�U�;�x��<\�2��
:�����Cc�����f�����Ph^�?c���=/Ӈ�E�A5dZ	<3we��]��t)�!5��r|�[�� 
�_t���.^Ä�V2����j�^+u����O���~Q��I�V�j�g�7|)�;<,���?jNr�b5�^���$����9���d��BU�o��ҋ��dC*<�z)�{�g��H�i ���֍[��
�H�1��U�]܈���l ��CP�6O�-M�[���]�����!�,�c�����A&]CX�vh��_mD�'�f3?�A!��"��T�nN?��V���N�K���He]ψR	������2����Pͨ�$�i	ı�Boy�Q��~`�pA��s�p&|Ȉ"�gHm�O����B٭
�����`ĘZ0 ��VGR��\��>��"�߳�H���g���{��=Lf��'�J���-�����<�@�����2�Ր��뙇}�n�Ή�=��̓�8՜C"�����
�	[	[�{>���"�w�-2���5l��J��|�Ps�g��@���*�֩ss����Ϙ���U��+8N}�{^U%Q�yq>H���xM�r��&��rB ��l���=��5���(N��72�o�3��ٙ�#R~�)w��
���������ζaQ���k�s�E�"��D��`�_��"��(�M����U.,���'� ̀b�������{y�6��i�'���aMz��d$}�FRWv��(U�s��2�	�2=�� O;k~N��.v/HG�Ũ�hN��5S�
�Y@t�AV7� ���lU�;�!�k������<-��E)�� �iƘ���y6�͟o�H���	�nQx�&�wҒ���Rɿ�ɇ]~Z�a%�Fd�k�
sO��<�������=.�kl�;yK=۠��L��}9'��X*�8�T[�:���Ǩv�'^5ə�:�P��D�ǈ�o˖����ʸ����zJz���kͩ�˴�}ח�n����`�>_KIpZ[��9#"��J�F��ee�txϬ���*}#B/�[��L�SjI������L��������-��;���f&$
<�L<����������@X��BR�Ա{��64+��w~B�c���ԓnla�]���1�-�`g�Q�D�)tsJ6R�x3�%f9<�&��6�'�V4���� P�J��>��'r_��)�K�^�w�V����Cܠ��*#�ޔ������A�٧���Ʋ�1�y.����<�3>��Ԉ@U�Ǫ^e�wcZt!�^)���̆s3�����(�|WT�L�~0��$�'�P��13',kTy3��͡UKqe��՜��X����}ʱMp�qsCe�R���s���7���.}6�$s����y�t���(�Ɛ��P*��N�����gF+��Mޛ��ۑ�d#�%����h���2%�4����I�2�>d	����7"�	trk$���ኧy�"�����*9�3��u��H`�6R�MG�c^���܁pE��+W��P1VV[�E�a���}�
��Am�&_Y$�5�2��iE[Nj� *D�/}Cބ�7Jc,N���<�����M2����>�R�Vm�C���]��~�0{\C��x�����s��bR��L�}�G]~�
Oe���jjH{y��x�^� U������N�}�<
n���p�����
e��{qG��\ǩ��3f��#D��"����72C@m��Q]� =^:>�)�L�d��"z9��@|I�b��Ǡ�rH�e�"w��!�l;ZT��[c�ڷ�<Gv�4m�@����DY���i�ЬtG��]���΀��џ#k�,��Bl�r�J@�eWg��G���I�Xq�-^����w��&�����w�P��e� �w�	/+�z߇}Z��J驫�-p���g��U<}�Ue�_s�='(4%F���=�4�����ӄ�3��s�,�3��n����7�B`�D$�n�%�\���L�(�1wV
�_@�~]�#2P7?���O�-�6|��ֿ������p�[�uUU�?]]9	@Y?[9a45guv�"X�/C-'<wT�B�Aa={j�IOs����Pןb EF��j.X����}�I�X�5.���\�GQ����R��v�x��8���Z`4-cQc�ճll��ڨu��x �
9W41'[<����f���U@I�`S�IQ&���Ԓ��&��=���]��|d"�T�Xm��W��Q^�p~�����E/�^�=����9;�����y���2�Z��;���)p0��Q�nK�g���yga�7�6~�ԫN�}-999pj��#r�����q�d��G����#�۷�}�� ��p���O��jLN-3�,b����9j��jz+�v��1oe&M�`�o�e�'��*�N�]O���[��p��%ٙ��3��^���	�R�zn����BH='��~�@���~��ĩ��'�����t��e���^��D�K=d�S��>���,�5�aH�M����NE��`_4�e��L�P�4�Ȗ��k��&G_��Nņ�oH��\�=�&�I���Eڄ}�ѷፃ����8d"�C����{��e�V�Rt��ON�xi{�D*��P7�
1���9�� 3���K�P��ܝ穰 �
Y-?���3x�Ѻ�����7�IT@=�O��;�;�A*�KxÙ�}\�js���9�r�[���L�3���G����2}��E��������?Ɣ���k|��%�-�O�ZU�bp�8���k�I�yq�� =�-�����k����t�rX���-�yJ�2��l�C!H� ʕ���6�Tt
[���=�S9�S��i��>���T����o�e,߇�ډfkqe�BD���3��@)K8T(=\�a�>���a���c=��u�̞�{�_��`���H�2��o�ϵ��dr!_h(�7\%����_��r6�EMW��F�'��9�';�Y_Њ��ٶ:f4�t�֠T_#���t+�f�{�������/5&����,B������j�Ơ2of��d�Bj�,�fn�7�n��1�\��{k�~B�NNŮ�([R�4�s�Kgo5,ԯ�}��-Ɓ��#4�/�7��E)�fvvz���
�T�A��;Uа�]�_���W��\��^Byyy�ؑ��Y��S$��q�������zF�����+ԕ��rP�X�j�k���`~��<�I��_��\��iK,e�����0LXa�]�[$�D��\��h����}ؾ�Ƹ0�)!w?��6�%u~���F��?����W,�����j1�\^�q<�vp�aJ�iAaN��ѪYUR����`�ʻ���5]��!�s4	6o��g�"P��AB�tN h��h�4�FQ���0�|0�3�p��ƣ�0{�~_������U�i��R}(�ޏ1�n9��&q�ı�����K]X�sR�C^��!1�WLb���A	����F��S�Y{0Qi{��Jg	:Z�U��oy��ԉ�ޑ(b�"�%��������>��k�4���l��#c�d��r�V���.���y+����]}�_h�n�KE'�A=H}���<l���%�S�y�ա�&�K�"�J7�kn��y�ȥPŌ�t���o��_6��h���Y S�3��@��`�0�U���Q,�E ���O���x��g�Sl��l""%ޯZ���4������CP��L_w���BZ�.�Z����<ꡟ��[#!�W3�Ս�u X�dx�����a�{��H3��N�PIm��,:�N�X� /�o�_�ξ��hw�Q_"X�-odz�ש���0 �ga�a��<�t�,�\J��Zo��񵪈��-�eNk�$����ZbB��f��K�����d��1�w��C�u��_@Ҩ�	���)T�lEc�d$g��%c���<�m	Wx��.�����O5���U7�|xb'��<��y���0ʤ��#E�z	��װ4���rS'��s�4�Wݧ"�\��D&z��#�V���E�$߇�%��ME}�A���x�� �Ș�vXa��7��p�?*�� �z��X7���e��r�8�[��Ed�Pqb	����I'y��+*�K�N}N�5HOn2�<��|��}��0����C�$&Y����,l(Q��y*f�Ն�P��̟v���WҖO�� R�}���.:�l�%�ܶP��������]4z�|UIEu��?����ΝHYh�C��P��O\&�;V')xv��%�f{��m���M�t�H���,Ȭ�J�%�o'X���#��ny<�%\f�ƌ��q` �[;ڐ^��b�7
������YV`�]�@1pl���޸��m�Zj�e�P���>u��ct��JR�ƣ30��>H��-�2w����h�k7Ϩ�r_,�}��@9��[Af4
�7�D��������7������E�t%EO�T��Ͻ[�a�8��dOGݥB��<��?�f�/�&$͒ݷB!f�����+~Z���*S���?yE�3����W-
ص(�1��Pz�����_ !x�����{[��p�]T������iV�-m#��]j�Ӌg7��T�y.�g���'��!y��E|��N���� ��jE���k��ę`Q����q�,��M��v3���w�_�]��C����}z�{��]�d(w�܃�݃����V�~�ﰈ��u^й�u��0$r�}���o���[:%�`u�~�������Y4�S�
b�m�����8kp����x�����^l�6��^{
\��=j�¯��L��/���rw�>fP��㒺����"xb����գS�آT�KV���=U�ˮ��U�5�3��T����(Ӓ^�t�ъ�(�ɲ���%�4�_?�mZ0�$������$�O5���U�]E�����eM�6����Y*x=T�b�ra\u�v���.K�������*`%M3URP�~��b��������&rW�V�����e8a��T�斷D+�I�/�2x��un���$��v�ZF�^��r]����2WTǲ�@����7��zq}���H�01�,�~EIII�r�j��&���ƲI���yF�Pi�~Ը�,�cy��GK.�fQ�[�n9���B��+�J��C�/�|P�خ�O �+3�ތ'��8��)C�,�� %���϶�54:��1!`��m7%�fZ��i^	}������oV�]A�9J�l�EbF���jp��$I�����G] 39���suc̿`�B_ƻ|�rKO�������0 �N��C�4b�k��3;;;;��q����՘��+�^y䵐>ʩ��XU)ݮ��_�� '�7���D�\���1 ��#�V~`)��iLJ0���m4�X3!�8K
��G�xF139���"�h� a�V��:�ڕ�m�*s�֚?�V��ݾ�?>2�@���I|�:*5|m�mT�����.Z<��k羄�<>���I��\�N&��au��(#ߊ�S��d��n�ܕ-������
��7��u�w���`<���F[i�|e�U�{��H���;|����N�x�=�&{��2�
�L����DUs�~�Pz(���=�K�_u�����o�t��I����CUF����J3�I�N@c���\]�y*ɦ*\��}d_�^��{ �-k��SkwG��C�^ޒVt�Ut�ؤ�6�*�sm���]hèW�Y�ӏZ�����`h�)�����׆g���Ӕ�4N�au�ȕ������p��ka�"ǔ��q��㖐mb��<i�78��:�E_F�Ph�Db~[?�;�N�U����ӧ#P�	�߿�џtL"*]�	�V٩�o"
�[;�m@�������"�� 5鼓���h��<l�Rt��<�}��UWP)@�7�m%x��ѕ���R0V������7¦�j!3�J��M�����G��=��@o�#�@�](�M'ݐ��tB|�Rp�Pts��q�{���r�r�xi�����@M���n�q;�۱z�}j6�����N�����o^������Z�3�M��˓[�Pް�X���*�2�q�y���511�L':�z���N�z�)�ژ��A�Lh̯�X����!חMK�!h�f2��'o�Ki���U78�wZ��!�9���x�
���I�R�O��S&#��a���5�Վ��n��^�Z���&��"�i���*��8�E�_qqqPs���`=��7V����/�� ���B��Ï���{�bf����6V!!eP��Y����jz#��Hy��p��V4���1�Sb���8Qʅon{D�ϯ�a�K��G�Uz���g���Ѐ_�i��J/w-��f2�6OT�:��Mh$����^/�5աzOQ��/t��9������Vw�q���S�D��2�7�P�����O���S*X�	�K��$罬U�h�F��u���L�a(E0o�ʦ�h��ŏ�ϼ_,���U6������Q�� ��Dn\�K�nha��]�H|M���2�tY{����!h����kY:�ae�q�'�B�����:]3�^�.���i�W@}5>��#��������[�E���㽾Y�v��9�~TQu��ZP@�|��Ʃ>�U��
o%����500�8�ĉ���[��V^-�)�*j9�X�)b99J{r�W 4��M����A���
���,G��xF#K�\?�l�^�'��EX����ʄwB}A�@�y1-=���D�,�Ím���w�Ըuf��^ ��0��ݟ���!l�6��Ч��H�x��n���,�L���_O�s-S�[(��At	�ƫ���X�&{j5l��J��t�TI���>=��j7�v`*���l�[0f�G.�%9�l-J��K�����>M�&��AM������?%EQ�`R��� f��4@��c��N��+�'퓯V�akEkK�J�����F��"v~�)� 
���n��㾻!��n-���5r/7��z ���6o�a���8��q�|�ҏ��`��P|o�y�7N��mJ�?{UÖ��^��e��|��#P����
k��#X���˕k��M� v5��S��(0�I�M�z��%i���S��D2�W������-�����Y���N��ʂ�(ɚhM���S���U��N�:rE��r�O�����ȾIy-Ol�LJ����s�Oc�\7�^s�_P��A�W5&OM��r�ܠ�T�z9���g�w��hV~�Ȧ
�9���r��)"�oX\�r
O$s�Ûۘ�NfF�%*QWG)JQm&�t�CoI���!Z)�f���6K}��Է�G&ZL�w}�8㓒 JI�ɓ@��n���/(�O�r1R�s5�76�|��n��x��]d�����G��A�k�P�S�������
c�� N��H�A�{�34��_Zoj%����N[�Ua4+5CD7O�d+��9
�� BO�r�����l����g��?�P��s��o�	g��y���j�M=}m�^)fLk�F��r�!�r4]2��u�[��և�y���j�L�}�����v�EL���l7� �
��ff�>��59�c]�P�Ivc�
b�l��/�Uf�x_J�T���l��J_���9��v�>v�gJ�v�L������$Ұ����"=��r�v�$l�����g"}X�؝��g����1�������K@�Խ�$��eM�gM���Z �&���I���B+��L\m3TC���y�z;8�P#��_�-��Th�Kզ��^
�GQ3A~,����:��9�jA��ż����}[��,a��e������O��M	�9!p���|7V�r����J.����r�����U��S�r��Y����x:�t�sfQ�b��#��h2�������H��54��o��*��4d�= }�u��
[��{NZ�_��(ȘZ����m�<[���׶џ�
�-.ag��;�Q�1��G�d-�1F��(�_�l��X�Qv�%���;h�����Fd��4+*0��B^*��mՏ�T���3T�ZP��R<uN�K ��,)}�iR�0�i����J��[�y���5�����;�/���	��_����ݝ��(<<}�}���F�+G�;�c����� u���|������y+��X���r9��Nh�j�g`8�MnCrpxd�D8��j ��=�XI���3�����^ܗ�ĕT�g�tm �pj\w�YL��!hȦ��[�{Iy����*��(g�|	.!?�z8��;��؉c��$��?�������A�//�I�v���rs����.O�$�l����4cw��2��8qjL?�2��L�ݹ�ǍLl����|�'��$���e"<[�Q��Z|-/+-�%�1�(��m�$�kY�k����OEh�ym��0�B���R����N=�뉶�.��uƅi���p�9'�?��}oM��>q�fR������~|�EG8�r�ߦ�cY��t����Ih�}&��jP]��2��^_.��j>��K��6�+8~���q�(��uEf�a`)5r�<��QW�Cڒ �cTqq�� �FS��/vޓ�m��p�z� ����P#Ҫ[7"��w?�Xx��u�JA���h�t�)#6�
H���3�K��u�R����a�m�����D�U��ՙ�p �7>8��\��tK{J/a��4���_E�dP��=4rZ�Zt�1}����q��>� �!��!O�?#�o��O�V���0�G��e��l�yÂ��f�^�m���RFފ��ips)usD:h�+��T?�L��T\ou��ON���l��h�� }x�P݊��a|[���Fܬ�ɼ���J��y�����y&Dʖ}�2aS(釀-��M)�����xJ���ֹM�H���?Gh�7�c��O��"-�G��e�����=<�t!�p|LT|]A��۽�C�j�o��,�A��D��ā�-���@��>�э�'�V�(��=��#���R��W��m�K�x�j���~��l_�
�N깺s�睠]�`��l��>͢KG�+�_��m����.Ĩ�����{����)=mj�a��OB&����`&�;f֝��� o�NQ3B�c�|���[ ���	�����pO8�x���=;�$u������N� k����4�m�n/G�,��e��Up��Y�T��S�[_L�~���Sj���6�$�z�P����Dl0ەw����V�� ���h��Q"A��LPj?�4��?�4�F���3��c<�#�ſȀf� Vە%�"(~���2���nd[^f�P_�&�u)�jxA�],)W%�đ�d~���nM���NN��WM�=}���0�Dr
#oiݻ��C�Wj�\)��?�������6I�&�k��d��D���Ԅ����j6c��}�����o���!j��/�.1:�{�'X��1�<��3jC���ݔ��uErN=��r�[�ˡ�����Ę�5*Q�k@������O���*GBd3y��˲�>�΄��q��cPe*�]���0�-Ķ�P��[^���t��{f����^���m߭�KJ�d�.�+e���h]p0�5�({꣈V�ʓx�r�X�"Ů���K����hn�ո�vi+�vL�X�.K����'�d)��:�ޫ0�������?9dS��ɮ�tdD�讄�d���SVG����EQ�l99Ƒ��BV��d�C���]o���{<�'�^�k<���N��2�g~ӯh�qiNx��R�g$��>��$��37�#XMuIa�M}�Y�^mB���Yy�~K�ːӔ��?� x��,Z���{�XjA3u��ro���{���F�T��(�<�m��}���i+?���:����n���k�v���B�����0���o�,��B��`�=-�;v��ș�e��m^���-�Њ߶�z���jAȟ1���c�OoN��� �i�q3_e�0q��L���ֲ:��%���������},@�z���%|�gpp�kx8k�+A�4Aڠ1Y'Nݼ�����=%<'*T(44t�m��Z�s�q&��	v�ƺ��p7JN��9 k�Ue%{(��� �t�Q=R�6������q�F���� ەo�ׯ��jjj�_}&�8��օ͗A���33-w9��'vT�~5U�q+mK�':��G;h��J��=��m��)^++ny^��M�����KZO0��s-n�ЃNyq�"K���_g��F
VPWW��q� ��03Lޓ��u�EԚ�u.W�Z
j��OS�Z�0�jLLX=nk}=8��u����2��������wɑ'^�|��e����=�%txE'�<�%�5���S5�����Ur���nCӱ�A~▽VXQ5q�0��sm'"x��˃�z�+����H��X�nl<���}a�޳ۥ��y��l|Rj��Kv���k�ќ�S��a~N��-}��:\37�X�#�)?=n�ٮ��p�F��+}�J��7&�i�􅋕Y�Ž�ѐzd�z%� 6��U��Ǧ��iȧ?�7���I���Sտ�C�9jUA˼{��j�%�Ec`_?u����@�7��"�h�!����'� ��$rL����#ZI�^����JW�N�a��4>8��W��A��'i���NL0ϖ����b�j97�e�b�L�����|о���(]"��S���p~��ku�]%%Ogg��С��̱�Dm��Pm7���{��W<�OM1��Jc^��$���ʲ�'��g����s�R�!����!�&�G��j^I��O���b*��ia��ӳ�f�%v_Yʟ��Y�Y�q��u��ͼ�b��]O�ۭ.s�6�555��v�h��\/��EEY
�m�`}G��'Y����72��yE��8m����=&��x� o.pM����P��ɦ��Bp:o���(]����w?@II��zr�I��tD���/)��+�}���}*�49Z���]���(��w������lV�`�A#%ޯx�����UE��N����Ӑv�=c��J���H��+�����D�Qć�⯛����C�I���J�x�z���>�V=X�#cxK��XS�
��3��RN��`���NE�U>�F�9�l�)֎%���Byu��*PVl��ȕϚ�z�h�c������'%����	�F�`?3���e�p�c���5�ϲ�z�x��2Tߨ(�>��������+?���k��S�E?Qǈ�V81���!9��z��v����z����ыd�2)j넄��L�g��h��
5��i"�o*d]b�N�!G�Dd_��x�	Ý�;����$m׭�	{�VZ^~�2F�� �|`&�yM�N�Q.4�^%_�F�7x�x\��/}��_Y��W��b.�[n��R���]��(��瘖�h�~/�w��g�=Ŏ����?��������,��OM��H���f�)���m�Ճ�|���Cᒔ�]�����6=+.Zb�G:�F��_#��. �C����x�f��9i��9]H1	��?�������1��=�> �PȞ�*IЗ	\H��{�cm+I���	)��'骺��UUn>�~qXwyk������������Fp�]�	i�r�Y��-�Я��x͟�������t�dW��qT�� �ɷ[�J+** ��~TĒ��K��7��D��Ԡ`kk�ãzb���`SsklD�[�34n��l���O���O=��l>��q����g+mi�d�jƏ
�>��u#�~���'�˴���@�ͪRc�=Z���������_�ml��,wz�E�`'C�&o�A��p3�f!�h����?`4^����'���iR�Q$ԭ����&v�+^ԫI�颉�Q�0r����>炶�	y����a��΃lD�)� �2�&�o1��2Ÿc�ֿښ}��(Q ,3��ۛi-�# G���)����Q�V���M��Y��Rl��v�==�Ū�K�A{=���0�*-t:���,U\.�H���a߉�J���"&/�Y�u8ꘙ`2%�?;��F۵�X(�,��t���QV\L�� ��W3h;��í��W��`�w�$�u����@Z^~S��9Y6��Ca������+L���f_�L�W�c{V���ܳ��&��

�֏����&�ߓ�X�������'�/����T�ѻ�G��f[��.'�/6 a����M���i��Vud�}a�;��&ݣ��зdt��|3��	�am,�%�P�=4����vS�o���ʰ��j���85a�@_��֦�&��m�ǩ����X��[iVb^�Q��
���hN@r\i��d�5�_�S������C3�����i}]+56�B��z/�k�]фl����OV�:��\5a���ړ��l��0��0�B�0�_JyM�@�qz%=�JF����vpx1��E��s�F�qvmD&P(7$��R�	h==K��~S�Ԫ�m�f� ���J�9,�����_���S���vW�R��׫5�$e�t���񲲱au2���?X���$�<_����h7^O96�42RN�iS� �D��3D�K#n�f��0�[����ֱ����wA����y��>�'����#0��$�������r<q*�>�2�GX�M�/n�>0O=-gQ�}�ڵk���Wն	@�$��Ss��2^��f�[bp�*5�F6vr.���e��<�u�H֒	���f����e��Q����TK�09�<7�^x���ԯ�ȫ���	�_����6~�Hz+���A`;6":�7��8��e�����YZ���[֨y�r�~��o/a��U(�O�y��7�ۏr#oHE��Q��6喅97A���k�N�@<��i���8b�_�����F���>" S�K�G����/��<�8s�!$�Ԉ��#2�~���;��ȾT(��i���+�#�0�T�2;q+`�����ܜh��r|��4�?؀%b��$tv�$&�͘���uԛ���ܸ}�v��[b��|&,
���Q�|��sk�7����2�?�йq����ʕ��6"a8fO���E��.���F(6���j(;�f�$n���aᎵ]yU�b�L}�-��,�Аkn����"��+�.��*��u���3�U��?�ؚ�32p�[��r���b>��R&�<Y�P��G��[�O#r��J7�^�3�pJ�/Mоw��%EE�����͟{~�2͟���6X�+��)��nl�Xm��E����j��K�h�dLFj%j�4��������13ށ�`��`����"%����҇;&�Px�_��V�?x-����W�� =rn����NQ�A�}	���aGBr97ʁئ�A_Y��iKȐTza����Ċ{�l k�*nO)�����a8nLHz��-�]^�vw�F�tPj�r��۰I> Zzꑍ����!lp�V9��*�؍� ) ��z頋�N=>�U�8]t�od�sq`�ݲ��7u�����;_k^	l�,��˃�tuoFV; q@��p7Z�����l>��>���0^�U1 }v�W[�s"Ƿo����w�`�����f���l��ӣ��1��	nA;V�nx�R5x7�������ܬ2ʽ �5�Ǽj��dۻ�a+�U/�C���Wf�Kʦ��I��N�e�=Ы�֏�.��>'}�Nl�A q����θ��&�B�w_�	W�"ޡ,&���|� �bs���gI�߸0P��R���&V&�c__@Ӡ�+9p���0��+�?N��S�������2C�ih�ӑ#l�7�n����c@������� 2��v1��Er�S"��%�
h"3��5��y纴��L(�O�ssHC�w���2�?�;dWZ��ðy�d`���%4D/��#�3(�)�%��M(]@U��]/����X�xAB[�kVV?�5�Q���b����
�
ac���4��I��Nzaha暎A��IX˱��}b�6�z��qn�0��<7��4.��H��0�}D=��R��7�
�^ �U,�=�m�m���������K���OT�Q[�k{�5�qP^Y���-u�[.�F������[in��Y6q�zdfhtD�����SH�_g�7�,�gJI�/^�|5&�`�����Lk{���_�0�2i��eI�vl���tU�GIc~�`O�Y�����p6@E�C�����C�S�]p����(`v�H���jLM���N�iY":��s���3a��i��_=�*�7\\��Ҷ���,��#������I�9Ɩw��l�VSgN���?�z�87D9�#]#�g3�e�+��B5���^l����n�_��X��f&���ي�o"N�e��0�����8$��}��y�Y�d��=,��e���vb̍�0�S^K`eR�\�~o���F��9�g�B�#�pz��<񔀂"P���~j19-�P74�n$�^�\�s�����--iZV�AbY-�4~3b7.z(s���ׁ:���+�R3`'X�ĚFG_������/;��4��ɖV��Y�6��ne�V%8��C���[W��ސ�X��T�&gg�� M��TVT|ו#P�"�N�ƕs>�%��Y L+)YH-���T�i��X�\��ȥqeA.b��n��E&nE�1�K�[�Xoؤy�X��jKQx1��NSS+(��ƹ��v��S}��n����RPRB/��J���t^��x�����Ye��Ҕ=}�^��ުl�(��NVfwK���@�z$.T(Џ�a���>(���uh1'�2_tm��P?������/<3��}�Fh@}ϕ�������Ձ=��:;��OҊ���I�
3g�1UW����8K�89����]���L\����|Lo}8(&�}c Ia��*.����n��u�R����vjMxhh:�QA�u�����{�P!&��5�vևրQ=|������xs �� 5��k�}O����Tu����S����ӫ��t	� w�t�t�[5��{3�ޚjSc�P��E�2��΍)��f�Wi�!�ӏS�l�cx����_�ul��O����?[ݍڞ�db���T�G�G���Ɪ��w��vWߍ��H�s{e�s�$drf�z`��u^I���j�;��bb���������7��45e�Z;#(���K�f�����{�c��#�/��ޮ�P���%��ƲR���V�(�����y3֜��s��H�Ϯ�n�d�92�_�~��s�'Q��G�[g��ԋio��{j����˳��:1�̙�-��d�v)���f�-�WJ
����:iђ`����tǽ�ິ�Sd��U�����2H��M���1P��Ir�SiZ���r��r���ai��#�j{%���Q�t���Co�H<}Z��6<��vW���,*�>x��2!�������C�+���;�m�˹���6�B�߮q�m�j^+'�g[����/�z��@N,M3�QO�Ac��>/"4�p\��p���"���~0�c�W��cg~�LVĆn��\�^��Z��9���ڍ�g�Oas|
����Yp<�A�9>Å�&�{�c�gN��h�~p3�����+=�a���̓;����a4����z�7Htwt!{����{�]n��F������kc��Z��c^ ��\ �1lm��C��\�	��k�=��`i��~*�T��5�Lpx�F��V��5J�p��\��\8��=8�}DP��(XN"}�:��6������Lq�e���r)Z�z�}�=u!΁���J�|~��ծ�����F_d���w�P�2kl@�v�YE�N�E�Lp:�ʸ��6�x�?5׻]���U�+�~[��&�X|�i��JoyL�p����{�O\�(��XD����1���?��uߘ���.���%���KHye��}]��xYi�(����NǶ�R/�nd�|@3� 3�z�M����J�Z��9���H�0- )��S��4���O+9P<Ի��À:gA�O>v�����������L6+~j������'w!�c��W��C�7������\�N��0ڍl"�#O�f�CY����a���d����~T�q�vy^]�m*����Nݵ�"�jS�T�LM�lO�SeUϬ�/>M��ٺ�.��׵�m�������u�YW`���!��f�BBDGL��0�^���)'���k
��<!ٞ����D|E���u�&�|�%f)h#���[=��,���!%�e�`�{�Km��0��u�3g1�25f�1>���h�ދɛ��y�Wd���%ج;6�q/�:y�	�N������֝�(�c��{Fx]��x��N�lI�<���,�YZX!��n޻����U���cS��M������{*P����N	����v���(�a�W?t��9�Q��,���W�������9�GZ�m�KD�M���!�t�lRg�݆��<%Eˊ禧
��wK��/T�v��i���z�*�n/u�,�����;�Ζ���>�hi2B�_
�J�[���Қ���?\)�s�,�u��![>t�ݘ�.�1P�E7��Q���A4�לk��7B���<H�%w���A�-Iy��H L.��:�\�M,�l��)b�;nm�jH�wePÎb �Z�Y��@����ҳkՍ��������:o�]�M��e.��Y��	�B��5
7���'�m$9?��~]^&<?ϢQQ�J����Klu��8ۭ�xD�.A?�c�{�@��WF$7���m��Ŀ=��g�������rU0fĔ׵��*����8r����yv�gU���u�'����V	�a��\.�do�����<�V�|!$&�U&\��qA�W�^���忱x���!�����΋��a_U������v�'�\<1sJ}8|-'��Q��ߐ�2�))lA����v�_'E#kj�SQ�/�Gb?�x�4s�w�
R�eqrph�%��s�j��g�_Oˡ��+����7�x���Q����#���URY����C����{��ث1�X�-! :�n���SU�V����u^�Q�,LCj��M6�G[B�j������ݏ��h�x4������n��R.]�q4f��׍��3�,���fM7%rX�J��s%&�;��]��H��+)a�]�a�Ar��ʏd�zZ�f0;LEM���=�c����� +�Ia[��d�O�����<�4�&r�ˆ��x��Z{���$W��
��Vv��B��ͻ/9c�ٻ�����#�'i�8ɫ~�����JOǙj��E�'�����řN��N�`�>��ؑJ�b:�[��;0�Uֆ�84S!T��u�XVTR����k},*p+��S��s����n��Q[q��\+'Rj��@���>����g,�J�%�
�Ŝ35�t=M���,�e"M@Z��;�+hik$�l����l|։{|�}��`�o�joK�Ӯ>�wX9K����QN�$B���ѓ�a������[A?��b���2)���:�C^�%��	ti��W)�m4�J111^��GX￧J�Ȳv��>�T��AWW� 6J655a���|������z�nd�M?�R\�	�����?t�N��Y,..�y�pa�
�����5'�����3��� >o�)uzĞ����E��~���;�βݗ��Č܋�q��LfG*�>�	�����w������&-��%�,��P�?p����ń�W��K몧"Y��g{y��Ps8쐙KLa�7CCM�@ch�+�o��-lSB�u��F��m���w��YEf��K����I��?��\��k��_���۞&���/��������;n]��D��Ǽ��3��ǂ%�<��&@W@�U۱v�kR� 뎮�������#�H�� ��aq�Px��X,��' ��͏fCa���G��B�3��~�e��&�����.�w�p�W�a�XE��}'B��'�p΅��F�W<�ǣ��u�	��Ӵ,E�T�IK�|隋��չo6����GHK�r4�P_Nq��RMC��~`���}�����sU���fl�:��7���ފ#�+��N�
tH���C��|�B�GOlWW�ng�
> ����Ü���>�j��#�HDw)��k�FK���1�|å_1����iPc$%r��Ng��+�r�<��F">Kv&�E�$BS���jv<���N�	`A��-�kE�Va��b�[2�u��Qx��/�ѩmv����I?]���ƤB�,b/�\�bJ<r^Q�(������.��Gi����4������t�0�2]ӵ[�����6��n��������s��?3��!-�i�G�Q�3�D�۬|�7����0���Mi�[�Iy<�,�S$�O�F���	�9���LWV�d�-��[ ��GOZ`��w�4)�y�\7EHk%m�2;�=�ug}RZs䯳}+�程�
��C�7H�jl�J����X�'�Ѻ4'�LN�(�ܯC��/,77~��E#5D�~2����.�b��!�t�f��F	TUlJ�*��Sb�ώ���f�m�i�A�КNX�U�9���'�Ze�}�/e�BM�u�[�d�dj.wG�MԾ2��>/V�J8�K�������CZ�^[��*\$�#���3�ϩ\j��_)N���ש������WYe�8����k��Z�����NZ��V�������	I��6��v�L�]�C�v���S#��7���8�`x{[�;n� ��>�� 73c⦟�g'��Θ����X���S uY:\�&���iݫ����J���!��[���S����џ�_�u�����Ɗ��`Z���D8��	���1�[���ڽ�ne��0ioY(����.+�t��Sct��[���}ԅ�V��qa�X��{Vw��oUX�8�bX|�r�e.����y���n?M8|������V[��=�d,�ޯ+@��?1�,�s4M�A/��9s�4#���WEA!ܾU�A�r|����:����/�	{dʽ	�8���:��)�*�*��g�SS$�{@�c2=h���h�|���VR�B�0?���ز���wa����7>��<�.�6';"����a�\�m�n���OL:b6�0���lJ���5�����ޞqįD��6K�/l&D��)����:��0��~G�4���|t��m�w�g�.�B�;h�  96M�S4���cy�1��L���a��GG��CI8t�����FM�r:@9����wV�p����'�لL3�B��lӂ�5��I�Y^|���� �Č)�f�u�ߟ�̬�;���%+���)����9}�wy����0�`�9�9��F:�K5��zIfKb<Xq��H�٘���Y���q$�m�+�e�?9�Z̟�9�PB;k&��r<�CĆ��Ѝ��[�&�2��.�Z���;��`;�sO���7]~ͬ=�[X9Zמ9޺�(���)(`b�ګ�~�KryUPקE��!���1��I	��I����d�#�v�H�ॴ���"\��q�� *~=xS�:tb>�ku7�M���D�u��?c��[������>��A�1mZ�X~�-��5�Wt��8Q0�����ҷ��'�����?�H$)5_k�on(3��:�Ǩ�!��b�jo�-�3��u|~vl���mf��X�6���o�f��d��S�Ҟ9������l�Gi��oi� ����an�+j@Q���iH��zV]~�EN��B�Oݺ����cz�H�@��I�O,,K+x�{��"��ne	�����6�*8�+^ـ�S+9��$�ZgA�3�����J�.VR�v��9�.�R_R���R�A�uj��D��>F�TW7?���q%��o8e�1��}�G}e%:� <B���y�L`n������~�Q$�Uۇ�w�P@�Ը:ܩ�����(����J����aFc�!9Po[S�p���Bܖ�4ŕ{�1!/�+L�����Ջ�:q���V�T��&��&��g��U���ׄ����������g�u#S��*�@7)[�݀�~f�ObE��(��h��y;}4П��+��o�3s)6GA��������̄)�6�o�5ٞMVJ�\���(��)C-�:�U0T�����C��ּ{I⽫�_��4�jeE4�]��լT����?Q��	�����,�A,��K��v��1�$w�mEb��I,N'������ �K�"�{n�(7)�6�˃�z�LW�� ���&�_�đI)�o�M^?���O�%y���G���7���H׻)y�EIl�^���DM$Em�"��F��-2�n.��C{��&
>�~�b+od�*n-����;"H}���ov����g�Y�o&�y6�����q^��]F�U���w����V�1-A]�����S�+��y�xQ$�o@P jȼ����Q%���u�s�?]K?�t���Wc���w��[en7+��I�_�����R�V^!�쥙~/��4��&�t�:��j����IT��FEEř�t�}��QԷ�R���"{A�j=���-.IJ������1�Xh���Ť�E�1��ts8��5B`Y��g��k�x��6����y�����a��ȿPUP~G���n, ����y�� �"���8����qY��4]��P�����1�P6+��;��wZ+�O0�����"�z������;�F	���Z~E��!4�2�� ���*���T���FB%{a���ȣ���=DE�V��K�W_�k��_�mhOt�n���Uٴ���:��%��q%����@A�UnУ�
J�LX��K(�p# ���S�b�����Yϓ,���f�R��֊�W�n��:�/ũ�dBW~����	��Xz����.C���g��=p�(1Ff�f^�ҷо�/3k�AB�md ��2�E�Qи:�1��)��f����P�����\B=<�t��D�y�m��D�ʐMh���~�]�"�#���X�_�ޙ�E��N�ܮ��8��K�,.�`�%y)�25��|��e2GM�H�mB�c�=���Ր��(�f?M�<�s=���\���aQ�[����4�����Tf2&��<f)�7U���bl��4Ѝ�����f%�s㦦AȺ�P��_�M��d�߻����fe�C �y�y�%3�阇E�ܹ��;^ vOW�n�ΝD�MŠ�y��ʈ���� ���;fD=ۺ��W�OL����6x��X����ĝ�]�=���s��R�9K�/t���B�����:5|��:,_'=���Wt�ǭo;m�CN*~�	��3��F��T<�$�gӦ�Zs�ܫƙ�r٭4������t�F�jc�#Il?�t��@�2	�O��������\8ﴮ��焯��Z |��B�$-���1*�hE�A��W#8t3��3*�BV��9�ʰ���R?W���u�I����.~�3E/t�z��m�sj����!��Ԩyq�;h�'z�� *���a�����!��~Խ�67p؋�K��������.g�{�i���;�_ɱl�
^�e�ZS�4}%���dO=2� ��~LV���V~����5
�*V��4����=�&Dl�Ww8� <Q��$NͯP]���n�>��+`�>Jz�0/;�c�Fi�=ˉ�|�:hS�k8�R퓝jU0��l�J7��j���{�x�z��� 4ݜ�z���J9�s���*�����~�.V��������!)��A�1�O)t����Y���E���L�g4c��`�g�!��Ѣ��gZ�+-��6�d2�ئP&�W���ș�R̬R�@�r7؆9eĺ�	�M&����8 t�nj�
�0K	~ڦS�ș�ӧV�� �֟�ӾMIk��}���Y(�^��G�����Kn�X6~U �o�`�V�0�R�P;�k�A�<"h-��ͫm"ٴnJ���J\/����"T"�^�&���SV���M�z��Ȳ�&љJ&�Ն� g��B80���׶Wt1�G�g�^іm�AH����ٖ�u,T`�:7J�̖8&P�K�6~��*�;{c��NP`YSǯ*}�es�	Š��Y�cA�$����9��=*��J�����O`����~Z?=�j	�-έ���F���� +�J����mm�Y��
z�gP�8��KD�p����K�di :��)�_@�3��t���g��G��_K�S��R�]S��{<��&K9��ݐE��N����4p;��xb�21��Rڐ�6�W�U���ՠ��#�3R��0\���G��-q�B�1�[&�����*İ8 ��6(�|�a������1� �N,Z��ǹ�Z�-�S��=! _�w��q���V%��O�9�
��}�p�u������&��yqhP'�N�|c'f�4�D��������#G'�_k��D��cP���; ��ԑ��0�ʕ����rm/�Y(��oefV@=�zC�.p:To�Sf'�$��{�T�P橺���V�6�D�����xF�����H �Ǚ�4j@���ȫ�l0�����PasLI\
�`eflv����<k����_
r�0�艀44�˄k�>.Ëߟ�?��dҝ� %�j�i	���NZ����w��u��/w*��a�����g�݃��>��������/�0K�~�Y�Qk�^:�n�_\3G���XS ?�$Ǘ�2�Җ����ʹ��DGr�������?r�ey-:w��Ma���q�[�_[���ɑ�^~W�,�ѻH�1;�}`@s�m���p�� �-m�t(��\?��;�에�7���Q���f>�	\w.��t}��J�=-�E�L�����a _�:��������c ��u�����$'�N[t���<���E���Ō���=��ro7F�,0Q}�|���A�������~��v�w�a'bC�g�G���cxi	�y��s� �8�w�� b�	�?6}Jz�*H������T���lD��=@�PF6�ȩ	lQ��C�K�j��-����p;�u���H�b�gL�&(=��G�����0��D�: ��q�@�����=��#��GI�8�_q�Ys.�7���RE��h���:���_¡�q�SS�3�;п��}�Z:7`3�����(cr�[�@�f��/�����v��G�s}�����h����r`�(&Q��ɱ�a��0�@ >~����Y[k�]��%��.��%���',�-��/������A\�'�_����A�bͯ��J	J��<}_x�ȸ؉11T�i	6��dӼ
+����
|/*��{���/�aϷ�tT�s��%uQ��CKe`��W�G��|~�}��L���=�ؕ�N����׻o�|@�@���J�i޷�v9�7�ԅ@O�tr;
T�>|N�LE|�x���_��C�,�v��M�gdPHR�&�r	��.�{��ز����y�N�+=�N��8���_�S�ܰIwݿ o]�N�+cb�_�3v�Kڧ~�/�1{�`��Y�Nr���.ՇE�eڱЍ"��a}7���B����LX����.RP+_H�f�������N��2 �.�3��a�Q^ϛ�ĩ;���㥷���O�lTr
���rf�y�:I�ΘcȄK�
�S~�����> ;@m�	(��bJQo����w:�S��U�f"7����M���=��nS�X{�Ӆ��>�"��/��<��Z�;�q�����(�wcP�,���Q�An���I�*�l �P	����J0��=|�$��d�h���ǾZs��UA$}�ц��-y�p��(U�;/z�!��@��G�ʵ��2���r!��p����;����;�*&�Lu��2���U_�z�7��A�v-��L؛�6׀~}�*�3��AJ��,Ԋ�s*��c�AuN�f�����۸P՚
jc�j�3/�ʄ���I)�`�u�t�����"f/���2�D���8 N�������j`�r���Z�t���F��g�Kb�m fRϵiJ�!̎���~�p�7|-�M��b��L.�Fj���^�6uI��Zf�[�ָX���@�^Z���<}�U�Z�˪M�@#)8݆�8k���,��Y�|GNO1V`�]M�2�Db�ૺ`}�>hx��>k�Ʊt�-IC�Gq�N�$Г�Tgi'��a���� c�I/T���/���x��6��� �٩����m�BR�>�(3	��5���$�^6���w��D�ۑ'�0�����
�pERPyL�(�D�65���/C�$�j�
0���J)����߂�E־}y�R�,�KJiٿN�d�g���y��s�-!�����^}���r��`�[�1�e/���-��7VX��0v�{u9o��?z�?���8ٵYa�ͨf���p����ӆ�l~�(gmI�<��>��;
��+P�i���a44�,���U����Z�62Pu<1�|�i��-�;�/��R�@w���4�w��9^9�M���B�2�s��
�e 7Q��Q�U)w��� pF�`�����]�Z����� &4�ŗi�l��+K�F~�{y��C�-v��y̅iMx_�k+��BF�u�<�q�w.��o�=�@�U��갾Q�W�Q�8�2��7�g}���$�.R����U�����@$O��Z=mt^u�V��/o���+x�l"լ�wI3_�[�Wԣ�/���+_5}�D��C�$����▿��Of�(�u`#n�O��9��W���g4�)��2N���{*������X�J:�����(�d;�J����'^;z�K�1�~�� �Č��	��r2�' 4�c�$q(����#�^n���%�Bhjن�>�ϸW#��"i��c��������5J�kJ�5�(y�6-�f݃�W�cb���&��G��J�m�Gu�)����V߻:�=���v�%��#��6�KhK	� �C�u��85��u���{	_���ɨ���H�^�&]W�/�-=ŧҤ[l�f�:�i�N-f��GA~q�u����7�]i��I�*�K��M~q�^#5�t�������	�y5z �@� ���t)(�c�ێ���j�J�P�����oB[d#8LׯH�⻼�8{�I���yl��2˒��%E&�o�oK��t��ޮ~X�_z�8�|�d�6�Í��PW��1\��h�۵�漦���\�)����w�_�c�"���B�va:�� �2�W���';	�~͟����
5RE�dJ�����ZK+��`41EC�%ߺ��k_���^��1�D����!�G5�͑'`hs炠3�y�+l8۱��������[�/[v<�!k��Y���T9K�k���'Ǆ�x��J�d�8I$�NU�QA؇Jd��6�:6�����(�l���}��n�W�l�JVOݫS�n�Q8L�K�&ĔA{����|A��
�>k6�VLNq���*����x�#���b@9���*����i2������<}�mF�ة����U�'I��#+{�L�P4}�+�������268�)3��:(�-!U��^]RcC1�F��lƒu�$��N��A]�������D���W������S���BMw�/1��I�I�'h$�|:鏁�����G�[������@�O��~δ �Ҫ!g� �4�Q���~F��/��E�\�'�W�),���J�2�u|�Q�j<�����͜9:L7�)U��	����5��/��}�ⰾN���UL,u#�'n�g��g�[x�o�ˇg�m:�OPq��Ԗj�DY�����ӡ���� :�����q��
�r���0���[NP`�������"~J.w���)>�~�XpHeZI%Q>�F�%����~N��f�hx��S	��a��[��|0ܦ��0�|���c�1*B�?�XJS��,�/FJ��Q.bp��$�8=���h��i�oD�σ�$U�.  �W���b�� ��FZ��O�9�=
�sʸt{A�'	fy����O�����a;�&bX�{�-��~�#({e8̃J�!�r�P6;�@���aiQƜ�FxT�����v �dw N�}a�3�6���^����
���%���tM�8�6��b$  �I�V�9 �F%X@��E3�%������]�DY��J+T������S��_Q��1l]L�e���;�
Eנ���kDFj��d�/Ϡ��@��Ρ!!�n>_���	�r��5]�H��\�b�|�̢(�0X�S�s���F$�`2����{Jk�ʁ[6��V�zH�y�=��QP�!
� ɻ*��gb�-����-}�?�DGX�oc��
��F��P�W�o�h7�m	�e,�b�k��Ą�h<%�������ʶ�<Q`���Z"/�Տg�0^�{���a�s%���l�������Q�P�"�ߛ�R�
�լm��"y9A=�@xb��
�;ٶ��#�y��,?�r���lBS��f��9J;��.�k�埰_�yf��\��4�g=s%���
,�D�ԻJ���d��m�1N��k����k������;��~"��6��l��iD�}!�qE�����S��5�����V���ب�A��%���e񺯊�YK>��N����D�����B��(�14X���Y�i6����F��s%{.3ᚏ��������0�f�+0�~���:�9����D��\�#�R�?w,�j��l�P�/l����|� cA'ЦG�{U��X�Z!&=�^���\�,�WH�Ls;9��w�Dn��sC\��LH���Bw��T��5��H�4�J���r�+x*ܬ#dl�,�S�k!���_a��O��5�S�"}���vL�	r��ï�R�������P�ǳ���"�E�{��i0�A��=��`����U�59KT+�H� ��0Uf.��#3	�����]��F���P8���/��{����%���fC�ei�}ɾ�]c�¨�-%*#�d#!	E�6#K��}_~����^��ԕ�>���k��y�i,l�E��p�h�:�Qe5��4�Ԋ?ߞ�mw*�t����mM���DYfg_���d����O�u.�J���'r������bA�A�js���� �Ӏh5�SC+���ʟ���8���Φƫi>H�@1ʽ"Q|����k,,�`�$�� *�ߒ]i�ʿ�~J���S�м3 �YF�+'�����`RE����>���H�f��B� p�;��Bo�vwQ��K-x���92w6�Q �,P��u���K��A����i�)!��C�3!�:��+��nԠ���n��ݷ�?9�-!��;43m�s�V�.V�AJ�;�"����]������'��� ���n�*��#�S�M�@��Op�Kp@�ټg���nnZ�w���/���3xV,x�fyl�-��R�����L�$P.�*s;�{s�(�s_@o�b�����&\����}ޠj	{Z׿�ê�.`��w7��{l.��ć�,C��O��c"}80�aնH�@_���xm�A���|o;$Q���r�R����'�
��N���sq8I~p�P6I��,@D����7;)�^���r��u��y��Yz����Yi�awO=D�P0}\/G稙AV��VS[����n��J���]�*KMBI��9��LJ8]���<��31��CN��N<
�+@���Dۄ�|��+��m��7+���W$s��W�5WQ^�ʹ���A��7\���Hh���f�d��^V�qm��^~ {}����T�+jmQ�<��'����� W;^�	Oɾ�u���jw�m���1�p�!�+��#���Ns��'��;z�s���������%���K'��{zz S��P�K���"�7�i��q�ҽn�8%�7A:��M�j��!�:�;��*��e!SU�	\��o�9f���)���u�c��R�#3�oF� �8������@G���-�ꑀ(M.f����3$UB%!Y�C��|Dn�	f��j˭���왯�6��a��7L�DlAy^ڿr%�\.����|?���Jc��M<%^�m�^�ؼ
 �4)�a݂�FN}N����a��f�9h+=�ҕ�(��R��|>�*S����ࣰ�\�O�{W� j!� D��������]���SBJ���,?G�܄���'�ɒ�ơ+��ӫ�n2��������"獀�����ujN��>�ۍ�X�4�.To�м��r&�M��їV��*tQ���@�e$k�2��Ea�j
P�q��y_����X�{-f0��c�����x	��ᖼ�eEM�BJg��!���֗i�� �~�$�R;���=����'?���
�>�����|�j�Z��.Q�D��R}Z�͖'?��>�,e��&
�+˛v���)n]�]-�����D$'z���y?<_x��C�X��]HyEj�2�,�`6�7��mM�����d��
�e�4���ܦG�o
�=x��r�	��TN������#��@=�r]L�>/���X��隇���,�QdzUϸ��e��@ ���������u!��h]�0���"��	J�zru�^:)J����|�f4�g���ɺ��W��,`�⽻Pc��NA=1��ح�����'g�O�@r�T��?���F�?�~�@�b�=�T�6DKL~�Y������5��� �F�ų'�e���ϟ!F�=�T���P�:���{"��|̃i>j�Rb��m�}Qjʗͫ�P �
�J ��v0��2r���;��r[bZ�@�e��ua�.�ToQ���D�l�Őc0t����jPҋ���&�d���!�H9he/��`f�s��>�8�/�,��?m�FhO��D	��v�����dʔyv�/�X��La��k���_K$�RV��x�IYEW_u���.[Z���Q�3^R�$��]=�=�҃`?���̾��3G���P�;/��f�(fiN�?SW�%N �j�����^�d_�5F�1�Rs G���S����9>����,���y<S�QKՋ��yM�FMsy�;'��#]3�7;{�u]�:��3_H��'%�k�\�t9�����RF {Ӹ#P. �xx�n��Y�e�
�~�,F:"LQJtCG���������ј��D!i�ٞ���:�&�܉.}!�w�>�>���.cn���ׁK����_O�l��o7���X*���8��%���mW��,� s�.��<�n\r%Jϯ�"�hJBQY�l�B
���t���)8V���f���ḻ���{���C{UlMG�M�i���}G�y�)��0�a1U�Y+�ޠ1�б�RA�fd��i8�G��1䘃��7w��i9j�dQ6��aє۟��N;v��?���Fy7�	���Ʒ���E�;v�z�����;n������x�K����--d��	,~��,�g���/�%TO�&9��oe��G�I�i7n.�p�wd��AJq!3���S�6tU�M���hzb����azQ� �7'$���r��qE��џ�����},�e���[�t?# ���W^QS�s:yV)������l��S�Y&��^�Z�7�hXIY�X��u�"��J�P_
n����#�x���'��sTr+������8HE�9�|�5b��$@8/er1c��(��|�qIk���ZW���J�$O�h懓�8iYI��+,m���o�/N�@$u{)��X(�p�b]Z�CG�cs�m��J.[Bx�?��"ק@1����KԈv(���XQ�P�^�W��ϻ��5(��B�Y����i$���E0�����g�*<�EVY�Wϳ�sS�_��3::zT�^#�ǦɅb�;�QjX��%���Qa�D���G���cJ�TF�^���d:�I��P�>�u��̈��U�@��p�෼G�ۅ�P����x��z?�9�2-���T����G�
���b��ʖ��B�k���v����}�@|<Aj|��	��N�s�r+�1z'a���"���m�m���"Z}�&;R ^�� ���B��Š"�s<[�tb��^�B� �>^)=�C䝛� s��p�2Rͫ�i�BT]���xux<HP50�ve�q�%mM[�W�^�Sٽ���h��E	Q�Ά_�ۛ�쫺��L�$�Oz�a��]�y�OInM���L��:{�*7��Ř�㣡0@�����R� a�8�:����])����"YV�f�Q:)0�!����OC;�dG�\J:+U�q�����(�[e���ӣv�!RS[�~��l�K��/$�u�����$$^��(�$�vx����♸�>L��:;��5��p���>����Dw{�I�  aW�e\q��xa+�O�?DKЖ[��l�������-����3�u4��)%��ב-[>�Ŀ��լ���x@6YmM^�fg����ϥ�����_K��d�ypZ�Dqril����j�Q�B��ӊ_��/�typ �2���Ж:�a�:�'0�N}��D�$����c�=�����b����D�6m�Mhj���Y(Q���p�)P }±�7�u�ӗ�5�5�*���X��a�x��h�ۯ�_���%C�Pt����`�"�:E�Ly�跂��"S^�s����͗�	�X�#9H�w(E���ZJ"r�"�F��:�pV=���n
"ݬjN��w���T#��6�8��ٰ��G�K!j��17]�9:�Z�
4��׮��Te�9��������wfbS���J��Xi��'�&n������֗�B�?�ٵ��J�N�'��� pv�j>��̸"��Y
gu��<�R�Ͳ6L('��a��%Y���T9���p�ҦH�O�e=�R�aQq�v�"Za�
���3�m嶘�A��k\��0eO�]b�NÔ���:vh?�e+Υ��i���|M>Ӈ��c��Ē��t�����>�,��q��ocϡ0��[������_��R������,�uf�pַ��|:A0��CA>����Vx�maz�	��x�MD�*H�p>�/����}V�٦X��\�VU����(FcVr�l2nK��@`?n�з6�r�4.d���%�j:�%tR�*ƥ~V�S��D+9�}���g0����{Z�6`�
u��BI<������EÛ��hnR2n�����8�&/C�b�H�(�Q�-����oiM�%T�ky=ۮq��(v@.^Ӥ�:}y �V��.?1���� 9���y�<'X������>���Ÿ��W%��h+�oj��2���ZC�N1[��2���¬� Lልo�U~�c7�h&�o�����B���L,��ن��ٺ���EZ�r�&�;$_��o�2�x�"����y�#�'�mRu�֎懎�@1�𙔺i�On�\�0{���LE/MݯHЍWc�K��
BZ�p���ᏼL���gwt�7��`
��;i��fώ�k��O�jbY
����-Yv�1$Yܐb2�
$H�4~��!O\^7������<ֽ�F�3am�K� D����>�;�ZPm���3�kotE�})>mQ�4nycn$�Q�vU(wh����VAg���?�1OJc
�A�=H;@�u��X�������=��SE�q�Iiۓ;���!�r�*��Ƴ�GM�����ulp�	 	_�4�(R6��(��ǎd@�����mb�U.|5�
mO��󖦚��J"ذ8F 2��z 1�b/b�ŧ���O?z�$$�Us�&{��}�B���ޭ�i\-�5a��s���)D�a���8��!��z��-K�<��-�W��#/�G\#oTbY�����F@��ý�w�8](��7�J0K�ݪ�w��3'{�)ϻ�`�K~��z�Qw��/�� �R4a�駜K{��5r��vM! Z+�p�������ӈM��*=�4�����&�O���:����?��{�������3��<V�Y	�����]Pi�����4�U�Ƈ�LZVtitF�XQ�d�x�`�
��)��<��z�	M�]E��� ��K�"�yA͠s�z����:�b̰���I�i��w�,�dU��j��F�Ϊ��`n7o��^��5�qO� I{��j�i<�F|��@�j{���o�Z_��d�H�Ķ�Y��������k\x�w����K��d�>+���.��vHz]�:�vO�B�H�2����S=*	�T0��3-u�v'����7n�qwY����$ z�ޫg�һ�ݨ)P�;���W�n ir��<u��kT�+��d!�b?<o�`ꗱ�T�p��{���|������E���oL��k��9�-o�hStyeA���LtƦ�P�j}��!/ͺ$-q_��c�IH�C`��i������	�)���iY�f%�����zfQ�F|Y��\FE`�[*��"�E�.�èB�g�2��b���'���cG���`��QBp��mH��>U��2Xp��ǯN�P��n#k��y �d[�3-�iJ:��"Y�4���˂a������g��=����*R����yr]���*Yy`�<`�`7{�� /Hy\�a�Ɵj�Ú�}ָ:Pt)��,�=��L�
?����z,y��gf�~�D5��oofy+1�3�yMӡ���%�Xn�z��ʚ��ˮbh���b�O3h��%^�Sq��	a ��=7(�x&6A�lT5���ٽI��ZBV���H�jͣ�Y�>��AQ \y�P�]���3S�������]��w�R�e�J��A����V?�:�5�rZ����|e�[lk[���q��iGܘ��'��;���2"���P��1����3ĳ@�>��k�,�\��pEk��ф�x q�4NKL��q�/�0)Ց��"�)������/�$�Y�ƴ^=A��z��U���z�}~�q]̡U��d�Y?�)��Hߺ���y({�8��n揤:�tB�_�(�L4$��<�O}�E��{mﯰ��`�y�vv��_Sϖ�`��1>[Z X����\�H�|,��k�'��y���!�6Jv�;�j�l�s-�7KI�XFv�
�u����h9���X�>�+Ϳ'@u�ɢ�UQ���Լ�[�H����#���J_
G�=�DH�]���i#,��k��q�h����gP��I�:��A�62<��&7���BI�Y���A�Vt�P#����bo6�	n�� 4��Q��B&��&������EK="2�W,�~N{����m�A�)R�����0��?�bM�@�|�2h0�o��\�ȑ�A6@oO�`����^��}�����u���w3�x4-b07��Ӝ���e#'�T��gu �*����Zg�_���O~ڐg�j��<�x�q�Ao�����y�j?0���Y�z+�{)8��,��x>(L ��@f>� �:qI./��q�a{�l�>D�:��O#T�P�df�nC�r�]��gI@�&NMv�@�F"q�F ��7~z�i�ɟ`P� �v�n�w;T���)�N�y����#-G��E`�o�+�` ̟�>{4����>�H9l]�A�C�l�&0���Wn�a��'�+�^��iG����F_�g'3����p0�v���j{�f���Q��I�P�i��*HxՒ��hc*����~b+��Q��P~�T���W�&��H`v�4VR7kuҨ`
��{����_gP����&�s��E�}>O=yȲH�4,=�@Q��O�f���������oщ��*#3a�{n�=�sh!;�x��_�C�"*�Ť,�w(Z�T�;�	�2�����oB��#,J��h57��֋�$?:=�F���y0��/T����l�D���"J���67�Hu�[�@�7Q���7��+i(��;r������W�;\4Ү?����CJ��)����jL^+#�v[C�Pfl2��5Pi>,/>�_���B ���R~۾B�p壻��iӸ��5����PR+kQS�n��/Fn�B����1}:��ӈ u/9�K}��?�L*�IB���Uw��Go$��^���̽#�0�ϒ���_l%�#A�g����E�:XaЀ�}��������k�g�r�Kg�VG��5|m�2x!��5��OR�=md:��{���%~�dkH��	�#��[���r�_�ڄD?����l�( 5p.$?�*9ѻ��Ч��Z�����>��veϋb�\v]0[����V��Í�5���=�20�bI13����=B��v�$ߡz������X��ca>���
�Pd?�N�3�u]�s���H�xZSo!��=g�vstz��E�����`�Am��@z3{GE���%h�FM���w�3��+�$<���{�:B���_���@ӡ����U#鏲�3�V�Ԕ�����2�&�r�&7����ѐ���3D}�}!*K[���Kʧ��#�m{6���7��3O�Z��kr��gO{���Q��, 
��y:�7P��Pc�+����45~p����mp�dme�5%[Ce�E�d �gbRa\U}D��bTN�j����R������8|������w�8�j�<[-ǹc7BYO��\�����A>��Z������k�f�\� �I2X���y��.w|�)<��S�������
��!0�E�������R�_��|�W'��� H�2��po�(��x]#/UFʩ��V�̹�"���^�+ Qn���>��{����R�)%�7�֯+X�#��Z0T�U��Y�}�S�"D��a��^$�k�E4�v��~g�у�bS��1���RL�Y��g�ٻ삉wv�0���<m����4�/K�9���J��R�8��94)����Ũ�cu{��~�ә��3���;s��\�%�^L�� ��bWP5��u�Fz
�ǒ�j`�d5U{�F�����O�zg����&�`�9�p�e���j�d�Z���1�cfӟ��p�o�2�>���)i�_�x���X� � ���$uzc\�)!9/F;�jEgqa��@3|�&x9Tvn��f�w�i���	�l����Ҟ�0�Oj���y�M��q���@����I�m~w���Ց'X=Ýf����Z����7�=,��tMѤ�C 9��5%�c���un�)�Fw��}>�����܆��w>���	�8Rd����d��Chq�<~Á@%�<<t��DX<�HI�#���5�>��$.��<ñx�[��龍l�Co:%���*���$ HF���?��Yޕ��K�����x��:L.����ЄL&��7�:�Of%�fM��2rT��@n��)���0
�Tm�����sj�����[#���26�����e�l��q�.G�e�Bȳb$��'
��Nу��n1i���ֺj.���X��$�� ��nsk6L�2��_� 8_h� ���:Y)v@��s��x�JX+ʳo111�v�^�@%�*5���3���p�c��_c���\W��5 qu��s~���'5�e�"��8Π�[�$9��/v�ߠ�ђpw$��H,Ҩ?�Q����ɺ+�>s} ƍ*��E���0ﱈVo�P5Hg���s�:��A�]�:���+f�gg�E�6/G���_��m9!EE�#��/"is^�{�sѶU��e��E��*G7��)`�@EձI�I&M9�(7OF2F�]̣������X�>���c�˾.<Q�[�L),�?d2{�isc��!������*�16�]k�P���̠�cpaq�hƟ6�jb�T���T �fy����f�Pԥ'?�~`nu����%�4��#&>������ЋP�u��X�M*qN�!q>���`��)�ښM��gE���Jg�m�ͫ%i'��p}����:knV��bO��Em%[��4n�+a����>=���H�nKG7�ڪL�h�C�5��o1���b�n�ׂ��TU�=��������(��
��%+�i+&��7��h�a�H�0k潻J{=='�[E7ި
�[X\W���.ǯ|�Ak
�Ǚ��4��������*@ӷ�$%G�$�b�ڜR�t��{�ڄ'
���!�W-@�O��S{���~Ku)D}�-;k�*�m�����Ru3BU�t�c��i���>��U�RCk���h6�w�;|[<�L˾a~sYJ$��P���6��բ�`}x�fS�V�y�Fk�`7+N�g������BN)r�p*� a�{D�����o@�]�172��#�5����z��#yy0U�C��vZ�c�,��*�є�l�ە���n�&�F^�_Zpc�G5�����^	���Y���ɫ�r����FX�)уg��b�ŅL�&r� ������D��H��
�O�H|�e5����WY��T�N�4�ą[a;����?������yE�1��H�Fצ�r���M KA��i˄Ռ\ڕ�Q6j���YR�Y�19��K���hf�b�NYm�Q��/-�����<�C:�iJ\�[H��FB��/�˓��4�����Z����bIQ����eY�Y嬀��<�Kk2 <`*���W�4����l��}~L�K�_Ɠ
]�v���of�#����C�P;5ۂ������u6�!>�?�(ٔ��>w����M��+b����V.�HJۮ��@5q����]�	��qǸ!P��P���[w��� 
��Y�F/�ا�����Z�>��_w���oi#��<{G��&��1)���u��]B�m��	ּ7#A*�-X�U7���V�9u5��y(4v�ă�C��v�\�,Ԕ� �c�W%c���
�-���Љ�3O����Z�|���v��fo.�����>�M�x���&�[y��f��S�M��.�����ZQқ���#5ɹ�Q.����-[��� a��Q��5��#�#@_��O��,=d�j=��'��oƺ��Q/\j�O� �{"�D�2����/��׃-�����Vb�7�pV�fv"
�-�ܑ�[���ZS��jҷ</7wGñ��2�Z_ RbN����cK-��t,-*�) �ӻg��jMv}R���J^=�]�ɔ8Z�d�
����\��R*�Z"7U+B���If�U�f�{c�C�{����Q���@��;��
T2�l���*T��]��a���ތ������JᑬPB@v�z2f�¼̆�R�м��V�}L��q�5��ٺ�F����<,[���E�=��	n�"ˡ"�������( �K��G��C�幥��m����"�����9!��|1ȑYf#��Li���*��<6�V��H}�Hӻ6mj-�§��jBl9�Yԉ��k8ܡ��ы4Us<_v�%đI���R�����AG��-LAY��V��zŭ�3\����þ�m$��{�����z�e:#�+4v�~��[�m��!��;'9� zp�΃����#;�e��U���c��uP��g	�LC5Q�-��]��jp�Wvg�I�U�9u��ï��z+5k�ut����1uu�půs2��^����DX��aUڼ�ld�鬧WҨaE �G��x��������TQ��1F��{H"���4���+�o�P�������/!�'�o-�Q�
M�FT~�}�y��sU���8��(f��`�."a[�t[j��������T5w8+i�U��]{4��Y��ƾ_vi���? z�u���׶��_���M�ҋE0��x�oN�/��>�� 7:����� ���׈p=l�����΀*g[+��(μ�.���7�:�N�s��}�����V�A\�֓��jd�pgVV�����a����=JCs��Q�sf0��Q��#Ì�?~%���+���3;���}<�����tM�cy����A<$	_��xgu�z�^�*TPϲ�Ok��&�l���>ͷQH���Y?�d��v�}r3܍Bh�>
��+i�/&��	��Z�<��\�?w�X]t([�8��`����Qlf�)�f�3�B��#ic������n�on�(7g�*�G;?<�whqGJ$Ǫ�qY
���<����N��)G��{׼{~D'+W�΀��
��󀟆ktu5im%��Wb�]-�۬�֟?��/%֓����Ê	� ���7���i���2�u�[P����j%Q5&;�J5�HJ�-<�a�|����'5��cr-]Gz�B�X����hX��!�A�7�%��H�J֥���c'p
����Tpb���M_�[!h`5�O�f�MF�]t����|���]���ӳ��c�K���z�^�~w�I'��K���c����J��):������Xz�	�����6!�?�M��6t�w��-3��I!v~�v2�s!x�/�+2�����3�g��i���%��;���W��"/ !Ժ����3Z\W�E g�w;6��bJƖ���O0q��T�jo/�!������Hn�j�+���/�V��k$���f��y ����<Kq�Y��.�j"����t��L2���4+S��|=jo������D���?t��N]?�V tZ���n���Y�&<\�|��'j�����4YYh�(|�3� x$��P�����
1J�x����qJ�FN�fH���rt�@�\>di+�A=�G�Z�_�x�_�UM���/��QI�� �;,�UVn�Jc?�l0/{�r��Y8kx�mt�Z�6�)�>�z��+H��M��S���}=sŲ�,]>�m�kkk��`��VW��y�Q��1��6��H"���	W/��hn6��ΐͥ�
|�.��,|�\K��z?���b���8W�ҶPp��U�������RH��\2�b'�����Wj���*�Ԉ`��Sx��������f��(.k��yb.d��尮��6�q*�,�yK�_HM;��K�qo�sߵ#��@��R�M#��Q�?�uҨ�����ed�Z��C���p�aYA{�m9��B�F�Q}����o�hը����'�����>�	��1�٥�JC�cXQۚ0��ѻ���x��T\�H�� oX��N����S��?%��UT*�㭕#�q�����jꜬ>n5��mO����Y5L�v�@êjj?&V�|ˬ�[�������1U.��q0�O~�Sᡭ��z<n�����`"�����t���gЈ����Ua!|�x^��7i����8>�,����y�vA9P@�z�׬$�j*�
��D�H�����&�~�l�|V��@�~㿄�[�`��O<�(�d�߲�Dv]F��P
��B��7�zX�,������a1K`
_�����4�u���N���ԝc���K}�,r���~u���p��,�}�e ��o]85;�Ĕ�"�@�K��bK�ɡ�죸�e���N�|�J�3n��r�`R�صnmc�iW688t�kCOO=[�u�2��p�x�K�؇��|\62Yl�O���0����]�fjʯ��󦿘`hX�~��G�p5�i4�]=�:��
������:F�^?�fNn�t�pIG"ǹ�>,vo����a��?>�[����5�PJ��Ћ\}S�����	FE��cZ�s�[(b:-lG��]�艠#��/񷜁9tX`,��?���>�4�i%Y� h> 1ZY��B1Mݥ��R��v:�8SR��F��Y�~0���mۨ`@>Z�ٙ�s�<񭭩�?�J��m� ���gve{]���i��ͼ߻������q)V�5�A���#l�}s��"�W�`��s��,l�;�c ����]�kdK�k�ǎ�.!�;���\�hX�8�/��6^^
�eg瞮�2���S���c�E�s��JM�KAHX��߰αc�ﾵ�{۴�&�jc��b]�Kɤ��9k�R>�$�k#���+����#M LJ�����ƞ����V8tc���A͖�>t�h����#Y����k�xl����v�w�����Y����ް��s����;��R��'[��䥜�k��X���/��r�]�ģ������^���`)�	�VA��Yֲ��׳
�߭z}��}/�bh��W�,y����VS��k�eD�����o�7[/,	A��n3�NO�9��ïBWy����G����Ѧ0<s��(P��Hp3��X�\��`�L���A��J����`%%H��-����|���]��[�粨ۃ��vL�<�1Ʒ�L�6��?̵W,��I)H�\7���<_���0\üԥ��ɝ�k�S�E�.p_۹V�t�C�΍}��#WC;��']W/pN�5 ��#�Շ&��cgd���`�7n��4�����4���>�
��i����v�y�<�]E�y�^�x���B��~���GT>k�cV�06�~j�s���ŴlP>�Ý;[Ŋ,��"�C�g�.{�~\ы�(�%01ݥ�T7���������ū+s�g��p,b�rҠ�����_	QF�{�1���&n��6�I1¸b��������, �f0��S�_S�&�:�1�;VwP��^�@�ha��C�q	9���t�������F�&���},��u�C�n²�R�t��OPY�U�U���K��;v�?TM2����y�Pw}������-������,¹	v�rɫ��)�@����K���^��i3Z��A��v3ͭ��}�C�o���k���k���4X���뫮#'���1W�5�x6�� ��ܼ�����˓m�e�PF�����z��ʍ$��7��KJ>-#��=��i�K�5���ԡ� `n��K���k��B7�K�KK0���b}��T}\��7�6��-c���pw���e�� �?Z<����5Pn#~|����vM~݌��gS�`�Y�8��\Mn�=gZ�aչ�RZV�T�D�#������7�x�0�F��wv���N}N|\�t�י)�o�w�9��cc�I�_���c���_���x��8u��6������^�S�98�"D�nQm�E:\���{i��|��O�^g�~)J�S��r�K!�=���S��m�K�8?[�G�/��:�E��`>����>0�� ~��A���L˟��T�>:#lI��D��l��ͺ�1��諔#e7F~<>Gx�-#~�Rד'4�R�:4F���̓�Ca�;C�^�~E<�2m1�����h'�Ӯ�T�o<�Ɠ�[�D?0`SU��Y�n�Qz~?���4c+*ԡ���A�ǃ�h�Ɠ������}�q�hR0t/%�!�������i@ּ�>;��}��V7+	��ƚ������w<,�����Kg64�a�`R��Y{S�������wR�'+�[�'�`��et��*-̍�咱�����?��D^�(V���v��3H�z��2�T8Rs|��"�:���ˁ�kg?�D����?����{���O�X�#89�M��Ժ��WU�G���T8��� <�+�,X�'��ݮ�[�+r�K�A|�N�>y �U{χ�Z��_�2�h���k0��O���/<aDS�U���������Z�lJ��ol͏�m�U���V��Vmɳ;�����pA��m��P�/j@:_�'so��g���54��H�ռ�F���nJ��<wO_�/Vgˠ�a��.��J�[2�ZY�l-�h ��
���V�
�32���T��$��M�w�G�`�z   �ݭ���f�7��&�qz���r��/6���я:򃞃�hk��g����NNm;J時�Nt��Rn����Ϳ�*�"7���"�"N�0��s�,�LG��V���/-ۨ&�'~>�;����R�Q��H{bIN���� �mG�f���*[�R�5�Z���K��i��!z��b+e��;o��x������$$��0�)t^���4��_��+-[z�5��VS�wW��ʑ���x]�;��2�@L�D�?R�����*e|yrg\E)�x��)��DV����������bP�p1�����U0�N�����q�̕���ʷ���0��G���F"Q��^7�a0�^@t���%��[�ԽN�<s��	kߨ�j�J���dM�S�����d"9�����Y*n m������l���Gg/��mZ�f�6|����N�p)hƥ���z���+V��~s�t�	02��h����FX(gŗ[��Ġ�Z����Ɇ���F�(+�H������I���/��e;JԘ�V}T�q{���(��e�g~\BO�6����(:�n�k6��e���99��}��.���Ҥ�%��[1�jo8 s�	�����f�ry-t'=P�H0����H��9u�,��IH��F��tcN�?j����*�������S��-��'�����3x~~~���у�(�8��0���z��;p�k)����D%}y�����}\}���T��E���h��#:�A��r�����UN��[R�}�x{�=���,,~N�@
�S�iwZX"�?][��$�u���ꕘ���u{�y��{��|N���X����qm}��Y7+r�UQ��QjX8�՘��{���5;6�`\�B#�`��T9$]�O��Q�LB�ԩ�T]x01>�vR@����UyI��P��O���o�
.�k�P4�}�E�eW��̬���77����wO��UG���h-�oW��X%�L��!P����{�5�^w庻%{;=���|}MF��7WLJ���:cW�|X�8����w�糪���]r���;��6�Ѽl)"o���,.Vy��P�z� I�2Q�E|aJ��rh�jGW�A�&q��.ǈ%��T�P��.�|x�g=%������^ڒ����lQ� O��m���%P҄,����||�XG�w8����<��\[��۲4-f��<���@�>��c��Ѷ�C#*t��$�O�w�6��]��K�ђ�s~�fW;q)3��>�C�Y�����A-�Ǜ�S��>V����j�9���
#N����&�d�n_�7��6|�$��;��*ka<�/� �g�D���ڏb�\�/`u�v>�O�15�����k��;v%� �c���{d�d�9���c�_H��6Qp�\���p��kx>X���5G�k4Nm�P`�E�Tt8�^��O|���ީE-,:<gHB�'5��Q$I�I��6&��O{��ׁK;0��$�ޒ��!�;�(�^kZ����Ky�Z��N�jhOn���J\�G0�!O5�����y!��������E�ꀢwS���&�o�>̓�17�l�_�[�](�
�"_�ʢ>��cϊ�C��À!�	zy��8c{\�"Y�,���#"����o���}�֒��+t%��H��o�4(��?K~G
��-@�?��rG�Z����P4=�'��ܰ ��û���`��Kp&�2Z�T����X*��-v����=-��
���g�'������䨰lה�)]�MN�K�"��A[�{��.�|����4C����b���%JTY[[j�>��S-�Z[�>V�b�18�=w6QA	,`?:�f�֯pm���#�+�.�FO7�Y����T�V��O����r�l���Ӱ��2�$l��.Շng�]|�z\�W�2K��?1=�[�BK���������:�quq�c6���ʨ��IByyC�wq���z@�wp�/ZIi��N���:���.SUE��Q?w��5:��\�����;Hh8:܃�HPsE	�o����]���_]}���I(��*J%��5P�ꕾ�:kk��JsZL�l��y�4WS,N��66p	��
MO�y�L�� ˶x��~=:�5:ܴ��h�vw�
��u��W�X�T��V����u@�W)��/=k��N�����TR:虓�P�i9������|�/�ˠ}�7�Ι��U`�1�&�����b�h{B����Q論�_��=q5�����Gj���*V�;e��ȹ��Ζ��dkZQx�oҴg����M�>������+� k�v��њ0cK����*�x������ǆ��{wq��w��s��4�ͥN��pxe��w8�k?������@�{ۓ	g4˻`�s(Ԇ@sҘ�\����l�>`0Z1x��������b]i��۴^�'����it�jV��\�rs`��\�Bu���m�	mL��f*��=7���[5s��]۵����i��������.q��)�ˎz(<��`h���P��O�o�s��'Iʰ�����w�ؽ���x@�ۤ�O�>ͷ\���wc ��2ld��?��S�˖�1 �?��W|��j�|h�m��^>.NʊU��W�0�v�ua�p���X忨�A�U��^c%�[��&�߅z1���xJ��9Ƹ�y�����RCS̴���V �߷����2��k�� e�tW���MgU�~�!Ei%��E���A��[���A�[$�F����F����=���χ��쳯k���{�;߫,�2����H۝5��7Z��Y�VF7��^�k���+�B��x҆O�R���LWr����IG���;,�Ŝ(�?,�Ṉ��~ޖbtr�}��󇏱��=�
{�ҲC y�Y���a�Kt�[��@?O^>$��x��\��V�����7���=ϳ���*�W@|H��zz'Wm��4��P������܌��|�Pd:a~�]v��M�VI��$���^s�i�X"58��xzz� M�	�����=�v�=��n?~�����C���q��/=�K_O����hr�s��}�B������U���59攢򭖓7��mc�f�m4L^j�-����j�jJ�8o}=1� ��wv6�g��c��G��|�e]��SD1H��y��V�H/x�bDc��t]ʿ3i5��vC���&T�y�C��5N �)��QI
��C���DY����@�o3ޥi�$�/^���4����z1@��V2���jb���i���������i�/��ތִ��̧�s��ܾJ��#,
�I��n�9�����2 ]ѿ�Ж�߈����G.��x&�j������ROk���6ZVx�#�=� 7�:�&�*Z���)U���R��Lmd�]9ڢϑ��d�X?�z�e5��-����	��E�iY�z�����s��q�>ŬvY722G���k�+ú����:F�:�pd��p|����Aj;,���m�ڇ.g5�Jļ&K��0���v��H���V@5��T�J%B�"u������golile%'���ϥp�7��s���=��iY��8����#�p:���L"_�=C���s�^Q_�.�;~D�!�|LY���n��U�&�
�a�1��6��!]�ߙ/]'��hS�����������_Dy�5P`�j`����N�8X�UM�z"�{U�5�p�,8�.I�L��_���߿��q�Ve�EO�O�KT��&W��������x��'%�����K&���	�o��D��%k�>8v3@�pU�l��d�
L�LGߏsJ�k���<c��R���z�4����l����k�=O˟��.u��|�8|l_ڈӯ�bp����J����ݿ[�ؙ��ݥg��"+tm��k�m��A3��]l3��~.�����~~v�S,���~�8u�;\O�j��X?�	W�5$���o��S���~�V�����ݲ�m�2B���d.56iG�m�\e<�D/ � ?@v��
���K��g�E���R��i�}p���0}�7/�O�g�N�$���5�����Q���H��ʩ����_� |�]"NQ@�1�!y7�n�ka߀7�KN;��1-�G8Gd����!��罓���,�����\��X�br�#��!�N1�h��\�m��q'��&�A����g. ��LF2b%�%3_�F{�F��a�����v&� �V�tU���I��F�fy��6z�L���(���og��lZ��AC��0C��0�+�ZN�~�s�¬s=�_w��pR֕�d>S�t���nS�����}��`����4Q� vN�6\��.��"$VւcU	ls~�^��Ĩ�l�F����	�����C���y�s�?c��v�߯=����,+��s޴�<4~��N��B���iF������+S슊}���1�gנ�� e�UWg?���.r؎�-��������aݏ�$��wD�{z�+�:�+��d	���G����p�`�"ȼ���P���ʭ��䎳���AhX�o���kŻ:7�(��I�<H8��	�@;��w�`D�	y�i�Z�F2{ڤ�tv�O�Q��o��p3�Ou4c�w����1h��m%�k���������㜇�LbD�eC�����ȶ�b���XIp���������9Ek�߂Q%�����u�1V�}�����A�">Ԋ��]�l�G"�Ӡ� ~)�myo�9+P�~�!��Z�̴�n�X?~Nz�O��_�֥�S��ʡ�����+��7�|�ꑙ�rƌ�]�ٮ��}���߃�{qN��Jr��T�^Z�Bw^T�N/A}�L��:/��X{��0�q�;�����������
2���:����T�ɬ�J�\z�0E����w��\]�a1�E,�C�62���Svk����d/�7i!��B���ʎ�<k5.}�?t;6��<�m���SL��5 ����;�:�G&��W�G�j�G`#����|��U��{^��TB��0)���&k�����mz$�N�Z�I�0hm�����AE��5�8x{�@�֝},Ϡ�R@�Kr����^���������I��sJ,��NayAԝ��Bqz2	?�� ɯ�B���e�t�ڿm�34Oɢ�P)q�Ęg]�0����u�ߧF��9��Wn�i��?��и���>֗�\���v�ױ1�������[��wd��ԟ�_~���s^"�ܷ�:an����{߸��K%:4̜kxo>�f�*S��t�g���1�(��b>�鿚*C�0sٺ.dG�丠]H�С{{�QXh��v����i�y���*�6����MC~��=�/B����.3�o8����&�c��2L�ֿ�Dd�6�`�4!+���jk� ������mqp�XG���*��}i�d�Bɑ���ς�����_c�h���dwW�-���Ps����e�|���'���P'��jV�>�'�6�C9}[��4$�1�9p,Aԫ��{7"�-�]4�I�Ƽ�B-��@��+8-2�����l�|Rd*�H��֥�L@u�á�#3�Mgݖ���_��T�JĦ���¢:��l��4�i]6~Ѻ:�����˟k޽�ʣ�8K�%~�}��;��Ct�|����#�VY�VxT��Uf�e-3ֿ`{)��2�#n�؆X�WV��5�>|�\�-=�0bՀ�ҞAQ�A�9�7ϧ�(�2���d�I���J���L��ǈ�<���l+?�QQ5���5JV���RS�aJ��{���VZ���[};ˠ-�b:c镊&���z,�0���\��ǣ�є�sYh��֛�����_����c䨬������R�>���۝벗�?h3�F���[+SŞ����rh���	��a�)H���I)x/��L���2�"?�A-6n��m��A���T	�2����Q�	��vދ�@�}���l�B�+7�w::+g[�չ��{k��i ��+�DC}�f��V�-��۫Ӏ1�|*?*!��sa��FP���3��U&�����`��&%e�mGr��[�m[+w���2����!��G�>k�t!$١H�����J��k�q��>,�W{ONk<<:zlD2�_�ONz<���Q�Eg�l�JsO�[MÎL%b��	�߰����b}WE�6�y��_ف#�� c�k7�qm�=���I�\�tG�[�����\l�����ȱ���f�V�S����!gக�Q[���)uЪ.��2f��9_�#i�^ tJ:LQ�_�z~�z�'-�=���vQ�a�xRXR^���	����shR�)�'kJ�Zs��l[�[�V]�B�1益q��f��Y���c'�.B�qK�q�����@�~��!��DEE��}^}
R>3�yCX��j �V$�;62|[�}�1^�N/C�dVOZn�;Z���lT�I�R�~�?௩YA=� ֨;b�T�΋:��V;$��a���x�j�c���k���p ��<A^�S0zCO���ο h�:�@�Fq懚�H򞪗7Q(���S�������T^j�>����D;�̊���b��0��Jl�������]><���ׯuUK�D��Aĝxhp��ߪ! tԉ}�+߻Rj��j0&�Zl��;]!��5���m��^�L?2���}rv�:U��3�Ώ?�t9�!2�Z��(\����c�Y7�uJ|�)�$cha��)n[�I@}�"9x�����4�}J���Ҳw� i�DD|�󞙆a�'%!q�A��Q/�G�1�sko�.�ϋ�v�C_��O��]H�tSUQ���nd�Sz/gm�Ĵ^�sl5������.'��塢$,�N�K���\rg�3��^ȝS���Qm�&[�$s7����7��p�8����JKqj�����I��b��󬵋T�l׋�n��7�^��%Ϭ7%��ht�Rʕg{{�|��|bb���s&*>�.N�b}���#Y81F�D��3<�)+�K4k\�ݴd��cK��-��ap��@%���Gy�� ������m@5����Z����-Ό�"��~�Y��c7D���ZG�x�W;c���ks%�ԖhE������D��"oCV���#y�V���C�B����a@��C(�CD$1\�c'Aȶ%7yu�'Χx$n�6��f��OF757˫��
�6�U��w���n�cm�u�v����-�J>�ɶ��[���蟲���s���C��H{��;���)�K�7��f�ұ��@-\j���a������D���p�����[����
*��ʸ��@�+rr}��t�b��z���Z�X��Y:��>�q�k���_����ҫ�fC!�'�ɯ��LfZ#��1q("Ex��� �tw~�Ŕtc` �4�T���o:cd=�9�Ix-������7�Lx���o众"�Lx��gT.wVt���i�o4�^f�����2�fY>�5Qri����O)3"aI�����!2�K��4��O�!9',�`�ۘ�B;>~(����W�Z��X��g�:����N�+=��	_('����u�_�r�����*�q0��j�N�l���L[M¸�Xdx!�W��i��X����1�xZD�T�}ڔt�����Z�a��['�#"zt9a�1����wO����_��������<`hQ��*q!�	�P�uz���A�	���(��W2��˱�DJ�9Jbz�6A6�.��7A�|i/�SK��$�/VV!M=��ڦ8��[��聳8��/�s�4nwW��f��A�X�l�GVm���<G�UC�`��"�1J䎜`��^������E������s�%r��݃�c������}*A����y��ᱵW�匛���8�=���M��[4�bB��O�f�v�ȸ��X����=LB���;�"E�<���M��Q��2��3K��,"Da���ת�p��.�����1�f}���TC�>:�uu9��s����2}������սo�0�#BEO�A��_/�
e๸�ʗ��S�a�ɜ�O8�VGA������X~������_��e��yWKF���a^�j��i����>��d�݇2An�&��6&/U�����7b��$�x�(�B]v։�tE&�z܄a��є%�fk��8P����M�{{/�S��z2%����u�mݙZ��9>��������!^�/�tGh$�;���W(nK:����4��cf���Ϩhu�����Zs�w߼����We&�$u9�{�~?��?�y�;(RvͻQ&���Ġ*��B2���T� ׼~R����CjF��DRa�1�����<� �C����.�v>�eOF�l��9rˤZ����1�eETux;������m}��[�y"��e,�j\4��HR�Ϙ3UV˕������7����FF*��?��,Ty��eX�6�ݹ���r�x�-^h���EK]��	{g�4�Xa��@
��`����g9��HG��\�рئ����w��CO �c����&��?���جY�t=�W&�m�����)Lm��\���2��^��Cȓ��w���BB �#C�m_�NLA|Iu�YmXK��z��e��o�[E���$%��0J#[�=�ga���z]_�:�N��S�K!�B��a3���MI(����o���}�����3�G�d%2�S���.9�/�T~Y$�$a�3x��HVL���Ցjn|���������ֽC3��҇�t9�LTP�4���J9'�:\��] ^��p�U�\�h)u��,�����5�"Gw��Y�cs��,y�W���SD�(�BW'��|�v�uǋ/&�}W &}_3=I��3ܖ���؃6�fe���V�Lk��_�@�a��Y�Ư致ȉ��������kyE���^�S�3a��>lz|�5Ж���]�������^̓fc����Ek�'��� ��G["��@�C�|����_kr�&aP��Eo�ŷc�q�[��;i���>46�H���RsW�<aէ\H��4��R���5��ūF����˹����끶���N20�>���s�����KA
�0���7�f_�`�	�z�Y����O
�?w�6 ��q� �~��}F��� 7�k�����Ŕ���Zc�~Ԝ�f[_z��tjH@8�]uo����V5����m���́~��y�&������w7TbOL�*y]x�=�'��SVl�U���ܸG��Q�I�,Y!]F�e\T��m8	���S呈/��^9�9[�1'��)A�Q�qDs���~p{���b�, ���RiȠ���؈:�=�3'��U���'�y���'|nO��r��7��,	yZk����ڟ���1�$;P��������~������"��PB��c^R)�إ�J0G��̰�5��x~�=�Z��+P���?�t���������K1%��Y���f[ķ�Kp{\����o�����7�4��y�H��^[h��\[uINX�w'���kC�ܩ�8Y����;�f>\V�wg_�F���)-�J�+Æ����iR�Kݟrn�~u�2/�������rg�L�k2ѳ�v��4�]�����������v7i�f���=�+Q�F�ë`�38�N�͠�r�e_��nM��\\\��7b�U� v�w�8�<5��zx�{wC	���2'�-�Q����o|M�r�s:"{�����M�v~CCCe�y�s�L� 1?��2l|����i���L���������A��2�����2��4�k��/����a,�F�����̣/���)c���]��^>M�t��Mܶ8�*���v�&=#���_w� 8bg5C&dR��������z8<�k��� �(n�hwo/gL�����8�o ��z�#����b[YY�06�͵�ѻ.�cS��=rZ�SY?��^	��&k4�\�斾��������H[��YC�@8j��=������:
f��s���U$/T@���lU%$L��Ю�&�%w�S	���a}�~BO�S�Тk��b�5gв~n`�Jab:���V��lsNG���ѯ��y<i
G��t��@�I#�4JxTh��+v�gg�+�KI�(���QS�^ۃZ����@!I�b�h������f}��3�1#iD�����\�:��8\�pBZ:�,V�d�v�����ڑ�}����2���Җ���t�O7��w��鶻6L�8�A�A���;�],`�~ΐJ��Pt����������i����^v �)f�y��(� �;��F�UL�ٷ^3����}o���	�(V��4wtT6�8aV�.��,���v��������Z��\Z�{e'���L*p�K��T4��(��b�������ƖS�� ��B���W��A�YBrZ~��Ď<{���)Vl�{�~���a���D�"�+m�s��n�@;��%��%?}��x�čLZ���I����&!^�L����O�XΧ���D������M#�/�
�IC��3~$�P��|��� K"��m�3ڶe6�8��[FȒ.�Mn�~�vsw���;�s9��O#�U0A.�c\Rw�/�!i�#�7�=���i�pp���Z@Kd ��4��4��gzi!�bg��u�9୞>�f*�˳q���U����mq@��q��	��?�fe)8KxKgQ�3k���鼃#})��	��-`���m]v�̤�d&}h^wy烑�ߔ�Y�Pa&I�23�-����wjl�)u��L����D������c�f��m�О��,�=M��47}!������=�=/'�������M�ƅ�Z��D+}�r�e�gq��
G�٨5��:��a-ψ>-nd(R$�|xI����=�Y?k�1�\27[��8P��_�����h�}�(;nB*� !���N�lh[c��O�U�q�I\-N^�V m#�DU�>�UD8۟�q��0�w�8���2J�����
�$�/���<�7s�6����N
�jJ�WNl-ez*.��y?l=��F�i�=�7Gtv���<�tWc�ت��--z���,yF)C�2�Ӂ����͊�@�$1?����A-`x!oѲ����8	��/jf�)�w�g���p!֞����ڡ>d��� 	*=
�}�!w��0x���:�_����+G��lEx��~M����egaꐉ��p<h������+�	ny%�n�0��w����l��Չ�[��q�
%ыϓ��+��J+I7�E�"�e9n��h*�o���>���e��f�����3��*F&��7�X��0mƴ"C%OD�"&	�'(Q�`�,�mN�ۭE�ׂ��ܹT� k=��ç��&^�`c�ڋ�Z�r�K�H�h��Z�1�RY���eR�!�3��k��v��j1˅�R����%/��)����6��Y�b�=��K���W�y��؜���$@n�;��iŇß��KoL�_��ˊ�?����7ܚ)HIKS�Ho>�BWS�^����쿇/N�'�<:}i�5W�~w�������]E �x��$+o⺝�F�Qpr͙��(�=��T��&�`������P#���uĞ=��d�1�����No������v�[��ZUX�~h�������k�� Ik����f��<�Т��9�k�����Z���t-	�dgA*��㬮4[z�� Ő�f.��k'g<���,�V}:$��B:yp&oǧ�V������VZ�h�8y=~��/qSաW����k��H-97��2vSʪ����{�v����CCٕ&	����SN ����k�,���l��WF?����1�N��Y���e��a�b"�)��O�Ɨo���������)���;	LH�1�+��A������BЎ}��b'�v]�>B�u�),�xI���l����㻻�oT�W'��э��yx�����f�J�h/}*�ׁ�����ɥ=�P�%�4��@LH��	��F�S2k�-o#1a�@1md���� q��OY�vF�_B
'@:�W"7�+���a����W��]O�ܞYܿ����z�ក�'>��;���!#�d�ћ(v`��X����%��!�Q-=������S�B7F���b_P	�`������&�x)T�����Q�QU�6��/�7�\^֎#��Z���h�\�=�1'q����.�<}A��s���;{D@U��:��əv��o����a<��i���S1]˯��H �X����+���KƊ�qc�I�Je�u��Z37=#�x���k�P����R�z�Ȥ%�Q�f����yᡛR���!G#��T4w��tD�?�������.o����/Þ�}�x�ě�&��{]E�a�Xt[fr:�Dq��eUf���.�����C"r݃��V���u�Qn��鴄�.����.�AZ���q�9� �i z�Oj����$�.YI'e�ǋ��ӝ_-�ɗ��}��	�l�Pd�}"/8�u|a�в�dZ���r<q'���n-S�z�'�����e۝k�~�ʹ][�������뉬�a;/��ƍΠ�PI;w��>ǭ��12c�q��J�^9,I��y�c;hׁF��OLW�����L�\���)sa��-��E
���]��7@�JY�ښ۰� <�1y�c�K�0�H <��h���t�7B��7U��n�Ϩ�@����i��0��g��N�>F��~�8��O=����I΁XnY ��.��\>κ�\�M�I�.��CM�e$8���g�=�"�7[bo�U���� �\�@k9��%�Ñ+�[6�&�{3Ҝ)�@�֎���`�����;}30���{x�sܨ��ҠQt�jta��&����cO:±'3���%���@O�s􆧐�p0��Oj���yX��F>��&c��'������E�0n!p,��+�qx����ȫ�D��\׭q����ߒ��-���ȱ�tp3:Q��o�!N���Z�Q�o�Z��Zp.Կ&�S�J��*�A����e��b����H^�r��Q3�8.S��A	Kb��?��y<��{�\W�D򒢓�h���g�' {�v+���=�ITa�����Q��&::А�뜂�2����O�+���z�Y'��Ǎ��G%�P̿�&�����2�u>�����{_��fs�'�ڮ�^�KT���?�ta��ׄBe��MD��%sJ�2���߶�ʖ��7�	ATJqqBC}�b�
{�BI_k��،�W�%�F���D���IO4na��7��9�Ҟ5�t�Q+.����"�W	!}#�gz0]A�X~䧉�`2���� �泀b�]E��qg�E�;��3K����P�l�%1G�n|u��)Y�>���B�-����{P�8��������Z{�n�VV��.�dJ1T�'�8(=�i�|Ϸ�cN48��CG�H�!*
�z,�u��L�u=!�����*�b��'��ɑ�]�.�&����*3�(�i�A%s{t�����uW�P�;�_��$
�HeM|��J2�TQ �?���ԕ�}��!��?�~�6�Ϸ5��x"���ɬ��!�if.Ш���I�����
?	˹�u�����`��t�Χ�Oy�c$uI�F76�@�oM����%Z���}��U�$44xҚ�(�Ç���zߝ��÷��`��LY^��ȳW��=|K���V�L�jFvw)������?.������+�������s�g��Xh��4�7�ōr9�� q���p�d�* Vh��kZ������Ϧ�y�P��76�ttj^�� U�6��a4�x~h��A�3)'��X�<	/c3�q���3�t둇�u��Mb�5\����X�6?�$*($47�+�9k����=w��6v��գduBB*����s_����7�G\�ZO�����z^7;�(�um]��7N�ַȔ�j�I�~w��!���~k<\��LR�j��F�O������'X�[`<U�1�8<G2�Ϩ�F���J	��
�]�5*	p�WKOW�R)���gԉu���6�hi��T�˕�����Ɇ�@oP@S���8�f&��8�Y
n�d������
}p�b����|̪~\��^0���$Y���cϕ0�����c�#M�Ӥ�E����`��Czq��������žag�����	|�g��s0�^�v�l�7����p$^���
�,9#<nJ��}i�a"}���0��ރOpٖ�L:�2T���	����h3��U��$kG\B�a \�{ X%�G6��mz�s�(@p<�|�X�; #�_z�����������i���H��ԭ-��<M��0.7�����FwLt���tt�e���JwkJ���m8���<�e��iK�����P����r=RB܎=�Ƃ�-C�ĻR
�C##,SNm}�'�[H�����/���%�xӸ�3e
-R�\V�:.�D�3*\U��B7aG�I/��\�h�8�0گ ^��aN�v�4(��qA\T�S�=�V�i�( P\��:�{_m>J����_��������Q��o皽n�y����o/�a�..S��KA
ϗ�I-0r�h �����~=Ka߿ĜB ��#�~�ׇ�.x�-�N�� �^�9�Ns�+&9��>�)/ %����.US���Z�xFt'Z{�/�Ʒ�)Q~\��z��XX{pl[?c���\Xw��dw$�~5�Tщ$�:F�w׻-����`��	À����qF~/���W).�P�c{������H	7���M,���!����f��]���P*�+/�����\8@/��m||�RR�c��vw��j0�((��<:��^ȴ�l���k����\Au�Ѣ�B�l~��A�e��]�ǐ(�ӏ\t�v��	�x���6k��$g(�VNZ��Q�v�X��s���<���1GϪ q\V\@�,�>���Q <�[!�����Jhn�`�B.z��h�D�d����: iI���~�/͍߅�X�v���6��;	t���M>)�տ�8�Q�)fG�8�ȝ���	7L��L����Y֥:L�$�f�jTd��ΪC�@2ɘr^A5>J	��5�&��|x�c�K=x�%h�ˎ��kGK����>��m����V�+}E'��[�{��.^�� �Z�?���)�����s�|pĹ�/�:�om������l|�BăD��t�N�勍�(�g�'����J2��0�F}�2��+�[��T�BȪ.�s�����0e���� y��~�4��%��i{/[EP��� %���6mq�.iDmGF>��0%^�2,gn�#������8E�`��ꚃ���Йw�4�̒m���T4�ޕ��++�BY������9����	�`�p�<�{���N�́�/��D��^�_ܑ7�s����Cʷ�ť�;�p]#I
��9��a����Ŀ��l�#D�Q�9�4K����&�Ƕ�r<�r�S��?!��{�{+?g�v���Q���E�~��Y�����R�"S@��('I�f��ﭽt3Y	�p1�C8dV���ez�6��o�E֎�<���0%��-z�*�[�N�]�d��^�.��f����u� ���r�����U�ڧ=�3!����zb��Ei:������U�L/,tV�z#� M��LA�-�]D/|Z��A���>�-�#3a���kw�CL�f[s5X��o��y�*K� }�͍��a�]'�����%�/޼�"CS�Y\��h���+���Γ�o�\]��\��wS5x@ 0圯�Lu�&�=�}+M��{p�X�%�p}C�vF�e�_Z�柗5Lӂ�7���U?Bڰ��� ���mIr��~J�������m(-��
��L�PZx)#�k�Ee�������nc�e޴��o|U Ot�/���'��N&lqNLL�Q����:uW��hc4��������i$�~�=\��v]~;��?tʃ'
�VA�@�����V�܆�l*��V:m�����$�]\����6�ŋW���>IR2�n�!]�^ihJZZ�Ėzhy��BJJ���)g�_~t�@O�Aoqz5�79H�H�n\@c��Ln;��[h�Q��B��N���6���A|����-�FX���d�g�^�����ǹ���@%F�B�O������i��N����;����WCC��	��f��2M<�|M:��)*gOo/�5��������^��{zF<��im�V+T\�	2��:�/�<��2����x���LgOV��aj��i���j��1/~�[xw���M��#�yFF*��}���i���y����X���~P硇� ϣΗ_����nȗ���Q9ݐ�����P*C���=#Ԝᖺ�b(��:� ti�rMٮ�y!�����w�ru�GA�%��݄�c �F��ͻ�º��� 
k��X~QE�}�˰'�I�\��¡�i*�J
�U5c?á�5*?�� T=KN�J����}N1O����ϟ�?,�ߟ����
^__�F����*-]-���5�M���z��jЈy��DsU�����+�������"L����6C;IC����m����5�PpGDX���(I�ۺ��%H6�3�,933��by�|������#t}�H�%�*K�y���`F�D� h�hTH�:�G�K4��ꭄi���5�4?�* �T�Lh^��0��[�ҥR��t��S�?6>zB �9Q�T?e��>@�GXn߬���G���ԫ�LpK䪘r
ss�BkcLz�^��c�E�W�U�W}��*�r��J�W*O���V�}_sxU���󦠚����	Um��@lg�)Q�i\֍�g�T�w�ݍ�/
�ۚ��G�ݬ��bG����j�A�h�W����#����~[n����d��#gf�S]�QrI f��M�ɧc�Q(��13�4���s&�M��0�پ������y��C�C������S�m��@(ɼm��Ӊ�rR������E�����h}�+�z�T��m����[H{��;���P������N?��_-�l�4!�e��t��>��q��U��ZGM���(qQ�V�H�`�_#)��!.M������x�[=|G��5�����uP? p���m�����v*}��a�L��"��w�>�� �C}�ɿ������DaKۥ�=r��t�W0���-{q��=^������kwᣟ�����������L��4�Ob/�6i����ml�Y|[}}aC(-A�Q�>3�9�&��OK��9�Xl^DNK�5�E����1;��k]&U堏_�ؽLt9�7�~��/uMp ��[�C%ȭd��]]���6Q9�~�����:'ЯAиD9��9S���� r�+yg��K�"����R��` ٛ�Y��`Λ�����o^�������3�s����V�>����|&�-�b[J��w�3�˗4���oj<�eDD���V��
���L0�T��'>=?�(%�YU55�2��YYY���$�9��b�rt��5�뺫ղ�(��C�ss��*ɼ�3��h�lC���[3N�e��m1Z�XR�����,m�Ķ�6�A��������8��˛�ƥ�>��$�`l�BB�8�⍥5�I��G9�Q6m�;]��Ћ'h��B���0�������ojg��K���y��n�0]V #�x�����<�j��l��A �=y�3�ѭ�Շ���ɷv�ߖ��hs���٤�����㪟�jl`���u���*;�=z�@���C���:g���FJ`����ŵ���8J����i1ql��-�פ���ؽP�?��m|��##�wԑ�	���������8^݊N�E�94���e1�58�7�G���o�y7j>IL��b��8���x'��g��!8Kz�[�����x4[�e|J� � 
fDO�D1Zp���^ ^��<���Я�?H�bv�1~_o���s�l�XiN�C8\h �\��!�k��hz�TL��v�㚆��X���1�ml�||��C��K+E�zi�*�	���t�>|�M�Љ�ؒ��b#�b[��qȸ�ԃ	R��#Y;?]�Ϭ���9���[�|S8�&_W>��S��o�wOހ��L�����ו��i뮦�l����DE�3��_V>K��Ƈ��e����%({su������t����(�r�2�����o�Zl��cFk��e�Fe2�Q����ݡ/���ޙ��6|�yi_��X�@J��6np� �1�!��0���w��J'�7?����FU�<�������;�����7oG�f&��'Q�n,�����܉��-�3�l#�,vv����32l���h�b�p��ٓʆZ54��e;��N�c���* t���YX��SD0@2w�U��"� �G�h�1 ]������\¸[��w����1�,���/�)�%�d��c��z
Y�J��͇�yK0���2v뭦h��
Z��la�%ȧ2����d�����@�lQ�ޕ}�Ճ��c�6�o?��\��]p$���\;�0��sj%f��gQ�䵵�]NM�ii+f���92��pdOw�Og&E��"BB±%n�.��Υ��Ƶ��~22z3�0���RԠk�@tSX�־�>1'E���/4j�e�I��D�)��w� �ƛ􍩫O�"_��1�ی�V"±��!ׯ�����z��£b|!�&�[�⯰P�o�'�v	�7Ϟ|o�̩��<?��v8����o�WA��c����&���a^���g��̦@��*�`�=R�~�Ƞ"��nC�������*|F^Z��D�B%�ϧ3�6��a��Sų�aq��PPRb�hw��]�������q/�Ȅ4���ޢ{�㰼*J ��77�/��+K��EKH�`��ԣ���>���_͇,����⢐\�$���̬:^P�|=�r�
���\�w:(<]Ōn����@���y��b7�;����L��2��t���䲶���-	��:���У���2������O�J^����ؘ��*�̳ܥ'�`=�r֓�M{U�ӟ$͐8�s�4�&��}��f�<�����	~���S�nA����qK, �g������ $�"�b.���3r�6��5�"Sh)�Q���x���&/�a�!͐�o�R�Mr����K��Z� 픬N���c���K�Ӆ�q���xC���g<"����̥�ޒ�[��S�9�s��,S�D�1>�2	}o¡� .�%G��{~9�r�n�3�hl���U�D�V�������E�$�-QC��H i�
?�4��4�Ӡ+K]�(ח�ڪ�'�崯Y�ig+��h��`���^�E�=sbUus�ȣ�:i�a�0�xv�ܞ$g�ɵ���fa��";{�:.Z{��9��4�Rє��Qe���%$�&\�;���~��^�s�o���8��&������Y���lL9�/y2�����!��
o�
n�����[��/�p�|���V��r}�ґ�Hʾ��hn�u���Wc׾��1�%}+9Z:r����⚠f����tvP�2yc� �k�'i��;f\�P�MZ�h��}��n�({o�A����vTK|�7]v���u�uB��u`���k}*ьP06AHLo`i� m�m�7��C�� ��3�2��Նy�^CfT�z���ң���wtFn��[��&���D,��4�'atfI1��u�QQ?a�_Z�I]$�n�%%$DBBZr		X�DJ@�KZbAJ�;�[Z���<�{�(�ߙ����\3�]W�E_�f��|���ȶD�\ ����n��]�n��Q�v��I���R���!��d������^8��cWQ��ǚ�2sxA����3�E�v��H�m�9+h
E�1i8m"�9v��		؞�Ab��;X��ڕ�CH���3�y�C� ӪB�c|<O����1���ߚ�c̴p�w�}Yo�JC�`j˙�c����1����y��L&�QaJϚ�p/��1���e�z���=}0��3'v�e��m/����R��ba��%��]���&��A��G%7��BE)\ ���ippmK��ԩW��#���ݨ�/w�w%(��}��$&z�Cu�d�{c�!E(�OZ�QK�(!&��a���c�<�oW9�$RTUk_6��̆�kTr�k)K^E+�?�9)����DT?E�*���vo|����R\�E�h̶wm�OZ� �D�Ҙ�;�r�D�!zC�	N��&�mrqޤq����[IK���Ӆv�|�&��As���p�
j�`��9��Հ�7��t�h��[���G�\R�9KMrJ?0찭(�0?���.��;�M ����;<��r&<��)����x�s��G�cy����{��N"�W�=�>CNL$O2c\"���Ӭw-�I:M�W�~�������H7��c���y=1�P���ƾ�g_��gT���d�>O�W�I�߱�O	X�9�� f���>��� �Uv�Pٚq���xWUc#��*���oݞ/_�v��������֯��J@�5�s���<��7o�r��EAFI AAHXX��tK��/�{��c�����'����N�>g{I��1e-�9��JKD]*C��<ٷw�Ҩ]?�|v�]&4��/�q)��%��F���D�Ndg_��Q�B(�͸v湔c��l�V �.,0�n�%�p��ؤO>SP�ǲ2�.��!��+e�� i(5777���ulfi9�~~P�}'����2L���M${�g����(��T.w�����
A�
�Y�v�_�N9���ۀ��۪�~m�"���Q�YO�S��8���k�q8��m<�zG�D�t{�2J&4��D����{���N�6�@ ds�}�B�ψ�♒��1!E{�>���P& ��)�2����Q���Ȯ�%+���4��r�6-�%�1��y?ŉ�2_�޲����h]�)/�X����8�n��(�7�	�wj��5�YJgfga���2�^߳�x@���R	�=��P^U�&�P��H	.]T��k�f����Ƨ`���'Kt�1�`�_�r�m^2d��ߋjW���Pr��w���o��nR�J��.�Z�0���l�F'�;i��Q�K�(�Z*��D���|,$j9􀗊�a�:WF��H�>&��QfJ�#I��H��F��咲�LN�	�4uC��K���%�3y���=c/���pv�5��Jv����@*0�����+�^�l����r�6�N�I���")Ca��/�&��l�p�;Gi�P�W�ء��ѧWZE��5�-l����V�?	�d�7:*�:��n�Z,}L'
`��~AшuRr�YQ�yΕ�$�4����aGk�x�Yb�<�6FsQ���L$��2US0��a���3�Ӕ]��;�|J���ҵ�11�6��ٞ�uU�:/?/���hD#t!��P鿻�[[v�Ҡ'z,��o��t�$V�u��j<�i5�hm�Í��}�ȧ��1�a�]�����C�E��S�����wp��ơ��.H��[yK�Bm_��@mc���mFA�G�ԣ���S��4.X��9��;\��/(e���k�|�~����$����m?�&������K++˷p߮�G����	X���߁����K'����^�Z�'���������%����&��h-�.��~��3�fŶ������E	�y��Ml�`YDI��0�"�I���=�c4��C ��Y��YrE�h�F����w���衪�ji�K
=HՈ���U���.Ԅ��E���Ⱥ-� �e���R�/[		:�~��b�A�h�}��y�Qe���e�Q�`�ޠA	jgJA� �6�3kM����p­��4E'R�&���������bP-OtD��z�̩q�V�\��17Q>�ΐ�_֔�]m�<򩴁�e����+�P��'>������A�U-c�goZ� L������ww}p�d`!�[f,}��G�"Zj���da=�e�K.�/VɅ
]��o545K��ZF��"�e��R��Jn��&|Z�$QkV2)�*�q
D m����DA�".����HH�Q_��5~���QC�u1�q�Ä�9�禦�Kt���U�P����v�gtyyZ�T�ޟ��百~�j�Pw�Au�9����R�`b�������S��L.��B4q[%!����[C�ެ�DV������a�� ������V��a�gZ�ӛ��wH�y{�����Eӷ���q�'Hě��C�-_�k���1z�T�3W
��!XwzS�eC��'Wwp�A�B���Ώ�ص,�媃��zlO>2I����U��W����H"��@Y�Pv�G.xsx� �&�e��qe����C��V��b��4�v2U��$6��fX�ǲ���G�j��S�}2FrF�������|�&��f�4�����]��$�{n���B$��b()�xDד�G�_&�5`�x�� MD0?�D�Pc]r������-�����±7�<���[Z3� �u����{=�����1�S3�,�E�N�"N"u��h�q�Jѡ�\8:x/�F�1>N~�2�T��Di��������d�O(8𿎅���!Q2����{;mÀ��'���-a��ꊞ̒��48�yg1�ț�B�G�}(Ѯ bMJ����Ev�Y�ŢuA$#��/����]����&eT�1x�ٷ�C��u���ͩ~2��sϹB<�윃�߄��������"�i����~�<<mX5�p���p1�N������St�!/��J�ҡ�y�B�ĵN������q��ׯ��ЛƀY(�gs%9茹���}���(�rI	[B�E��||��hA,V;��x����Ϧ�zy��I���5� �-��\Ӷ�A�_!��"d����<�HT+��I?%$�@����L7�@9�v�H-�8F�7+�0�
HJ�q"�Ǣ#r#���[�K�r��wα��[u���xR~��Y|�
��/��4^9;+�~�f+�U���ϒ���MX>�5������D��)�B�whg־gӿ��j����!�Z4���PoD  �.�%�.������㵷�P��9燤���倮��T����8������+�� �.���nynn����6x��*Lr��4���q�C��=��Ȕ�G�/$�+����pp��Eޣ�a�N�ϩ��ٸ*����~̐��"��=�it-�� [b�n�ǙP��es�3��A�[1���y�� ��n*�|I���\zx�=�7��sŊȧ�q�k�M/G�r�1AP��	p�؀��#�f��lC�|��&�g��cJ��kAI�Rܜam�k���t��+��췹��mx���y���H�����Ŭ	4����I+���ti����uw�^AUg�f�Ɔ�������*%���z���)&�<$y��;��a5Ů�i"`��6�p�۷�9&�߼y,8�}x���R����`�V�)@�{���q=�A�9����1~�Cf��3Kp?�lk�t���5���ݴt���ca��g�N��EK�D{�gr�4�Pw�A�L�)�M��D����7��5,>*d��9C$��� �\b�i9�P4��)�!???zgǝ��{Sn.9��#�����dƥvV����m��шU��	����v"���񼘥���T�V ��e�l>:q�X����������8;NU=�v����_z@8��H��B�
u<3C�!���)Sh��w���~�
�	����P5z�?�lY��~{�4�>�a'K��� e �ɩ)&g�啟Ɏ�s/�p�`1
�˷�9+H8:�T�����4���(̴�2�\��bm i]�{$a�GW��}p
��q����3D]�C�o�@�G�����H,�ǯ��sQ
kݱ�N������[�5��"�ìպE��[dq'|�A� ���N��-h�ꄾS�&��$;f{�O�����x��K<��:�~��	��"ɉ}_z�$�� d�@��L�R�����������@Xp�P�wꤪ"_� ��ީ��ʭ�ܡ���R����%)��u���� ��*�#w0��
m`P2 I�5�.d+./�sQ[�k(Zt�b'�m���f >&3�j��x���(��x�j��U��ü����0�qt��$A�ĹR�G �${�4WR}�Έ�gC-T?^����˺�p�|B;٨�vV��Le���>�z����Q�)��&v�����(�'�q�+�ٶ��߻ s��\)>	*�9���Ҿy
�#qO5�fgu�N/�@�2����h�JH��ZT2^!{fgi{�}p���!�pi���A� t���'��	��ǣ/�gR�@,���4Qמ��,7(����`	dc��W��x�,������6e��e$N/>��A�Y��g�B}���]N��
��;Ƹ�^�oǗ�?�[���\%Ʋ�O��y'��a*Ùm�FMNE�<������C��U�&�rƿ��T�(2PY�
�%�~��'�Y�5M={J'����'tx�Y�t~(���1�K��a���!M(�����ɿm�슺:�A�����yh	�h�J�}��E�@g�wS"��q2��1�~�������w�Vm��5:�<��wOMLA��:����}}�f����ڏ�1���QHzz_�`���)^%��-�}-�Gm{OcUa�<:�m~���ڿ-�_l���c�J�L�]�]���0��a�����͹��J�����_��y�?j�F3Kc���ҝ����=̿~���� �L���������ӽ���k��;���I0�f)9���=�P�B42�صG����u¡K�ّe%�,Mu}�u�\y�uC5 �����~D�mM�:`>�/��C2dga%'�h��C�h�T����H�5QL��Ԋ�3�,fh&�kFhH�Q�����|�`�JՔ"	aYB�!���e�NGO�(3�3��H��X���Ã����,�I/u(�H↕���L��;��Z<<W-@�u�o� #j>���q:َ�ۋ�s6�����ϙ�����{6u)�J�b��S/�<i�{"ԗ�2ד�gO�qN!3F�"�gͽ���H�A?�G���z������n�����X���7�f��;CI`��R$!&�}�#��5���,���|����ÿ}A��k��BܠB_K�]J�>���|�Ƅ��+�0����Ƣtܥc/��N���EO�HJJ"7p��=�&T7�0�� `V �Y���ȍ<�o��x������:ߠӜ����F�T�F֐u��Q�г���^
���B��+ߕ��~����6�����%��b�D�O��?<�:n��b_%�����,�da��4����A�2�?�D;�!�"�zN��l���w���e`����!��sX�ݺET�75eLYO]���j�ϩ��C�iF�r�y��Ą�ë*�� rRO�%�q��0���S�D�^^�G/�n�_�\"'�:��Ѻ�Ǒ�W�j��a�Z��c�_��r��Tw�74��چ���e 暰����E��0Gs󜃩���ة�Ci\��ӑ(�D)�q�Ũw�@�����=�;}�vƺ�/�#��LY=G�D;�G^w�տ��zT�2�E��^�Y=@�RlA�X�9m��Bv��mܴ6��^����G�΀�����zc;�_9�}�w�� R��Lsy3?�o���z���2��"����G���{�7�U��G��e�����GJ���7��˦�W�/O~��T<�������53�.�3�ݽ�?7�1�V;i`d�owo|2L�|�&ܮ�gX�5��aYM���]7������*-7� |���Mئ6�κ���Y�� ���������u;�a��n<�鹈0$����$��(#���yP,*&�ے�O$� �OD\\{Tm�VГ��!2&�n��f�)Υ8{e0�G���1��9���U�`]/���*4�Di��B��(=v_����DuX25�-�}~?�w.�*_�t�|���ҿ�^�dT�@[�4�â{#��bLp�0�#ͅ:F�6�2��v�,�@��t�w	�k�HS��_��*���v3�%���r���	fk{;!11���J�j2�e��a-)��<uH�����u�}��ʦY�L��Q>8rG�9�����go5ED��쐅"���So[W�܅$nm.��ٸ����4��w!3�Au�����.i����,:h�khK��z�� ��d��g�Tl���c�^����D������Z�.�A�7*���٩|aC����,3'�j	.��� ��O�SD��0�=E�^GS��=�G���eф�oOt��\��1�>����Ժ���6>>�/�)�x��o�S"���D�����q���G��_�����&&�n�F��NN���T����P�a���
���˓���j�C���J5�i]^F*i
�<֚�H��z+���<~t�\,d	~85�rU�[E�c�I#:�a\ҕ�^���w�S��"��n2���\�H_K.x����Ѯ�꘩uܿ�9x�9ã�1+��j��S|6o�ϲ�]N,��#�6������j5V�hooOQ����sk�TPޟ�rs�'��s���� Ǩ��&T[~t��[�w��[��;��N��4I&1���D�����TUUU�r�T���WL&���h�p2���^)�T����{~e���cCm���^��p�X��ؽc���Be}CP��Av,"U�Ґp�Q��'������j���6��C�Vv��d��f�Ys;�"���q��۹o|�ds�<�Tߥ���M�����6����\�y�9#6��u3�J_�i4�m՜٩�C�t�	\^C(�`z�l"RRq�D����;
���HC���%M�36rr�E%��� @����vya#�PZVF���3;��9�s��LU Cze����X�-l�v:������4�L�j��շj#�N�L�����k��2��X;Kxs0�m�]XmU�8������0�'� p����ё��津�/�f���yI{�qs�~�"���7"�ƾ�fe�t���w���s�@��8�8D�E����ͮ���!�-��$M=NHDt���٨fEM�����Tt��}��	�>'�XQ��N���2��@lni�`��M}p}�rE�g���h7;?��jJg�,2*Jy�1��T�z	�^ѝ� �Xni&S&h�*��^J��O ���J�&����\���r���#7��|Ȍ��w�����`��W�j������4ў���U.?��qV���f���r�O�3��^��g�F�����-�yo��E�j�2�|���Y�����뫢-�O�1G��0��xJ�4�]C�9�~^*�55š�q�4����!�8�\u�cz��N�s��@�pZ�� Z[Ǩp�Ow�1e@s�o��k���oY�-���0-7��ָeR䟷�O��lR��}���տ��j�#8a{|痥���z�21��������U	���/��X�D��"��1�� El��-\�B�����p[S1Z����:����M��DDj�%��p��(�*��X�_�tu)ߥ's��I��:���[2Sf\ƒ1@������Y������\�#@M//ԇg�^0f����9dM��xT_|�hf�9'����,�K�p�jX�ƀ�����h�5�tD p��V�ɟ�6ǲK}y�Z��튴P�=�\
�_�|����8N�ԌI�
Z	����}'P���O�p<����RDտ�l�s�_=�9��s�����ί�_��u'Ya��c�I�Kc�@��f�5�@�(��x0��@n(���E٢
�t�ڟ�Ϸ����-�m���PZ|�2f�^A���H�DH�\-�
}�T���o�){�sc�=�(S��mtV�@�YEAA�|�z��S�k�ȶPw!%֥��Ԗ?��^�F�X
�JH���
�!���rk�:�OL|�HR��ud���+2�y���Ge���&'��hL$��E�x��%ڊ�xE_� =�Ϸ��Iwpa��dnnn%��瑸8^b��be�8ii�QMǋ3#��h��xO^mb�����7�P�q"x�{!3���b��ͱc��2<Y���մ���ӻ��Z "����p��_� ž��-���}�֌,*��G��Qn����j#�u��ȕXy4�:�08��9�BL��#q7���)�@mt��zBh���89V��E�P�6�[�4g�kޡ����U�z�v\����%��j�7ul�ʇ�{�:NN�5K���_\x/��o7V�Q��#ub��Qb��e`�X_O*��ulfcs�q�i��ti�2�䕵���������d������3C�Q2yP�O����Ԃ[���s�٩;�*�0�G��������-�;dƜ��bn�d9 v�pg;���n��e�6R7�r}�'M�Z��"�VqIު�A|pi �X�ծ%dsj󌎮��c�TAO0��\��5��w��Y�n�$2���m��>\�-R9��s8U,�3�5x���lh�:�O��HJJ�E��Λ�N�MM5�Z�GA��J��r�m�}�������-,`��ᬭ��F�˝��.�ONO�TA�~��upV����-�y�a����=�+d�P c [�|�a��꺲�6��R�:C�$$����#��C	�� �OH޾v5���Y�Q��sE��ﯭ&�g���V(t������vS�0�(�f$ԌpPr.*+�~Ґ�s�����;9Ik�#E��~��
�S�"]�]ABd+��g�sk��)h����[��)J�aSS/l��5�fjˆ�(�����iiiI�u8_301=�D@c�He�������S�G�X���Y\�~J�Pg/��oQ�,ꖌ���u�R
��N[aDd&t^PAJUX6��(�� ��a-@>p�_{C���$�)�C� �����t��n��&�Ǻ�����	*���b���ʵ,�K�[Ā�lC^���=wuq!7.��Td�*�88�y)��f�����f�-l���!�n!�伀����o/�yh,-'��&dJ�������mG�T11�Q5G::���}�O2��!AXR�#06���	�O�x�H�_�EQ����Z�NVl�����]���u}C6��hQ�aD�tC�
ACk(KSk�-XN��P�X%8����ǖ��ƕ%D)d��ʶ
|�2�痒"�),`��E>n���&M6��y�!wWm����=T٨߽����(ё}�C��z����^��5��w,����F��^�
��s����j.
�J��D�٥�f�=&���!{���h�4�`��^���#V��.\��H�h��dB 2�V�'l)�i='���sm�� �5HK�4�@.oe`���m�o肧9��r�R��3�qK6�mŖL�;�����I�r�<˶Q�t���F�����*79HyUU���嘝��F�A�'��Wԥ��i�`9}kK�_E���$D3K��|gbb��$�;H�⑈"66��_�پ���"6ddd�}���� :7�)�	�diPto�+����<��2��;�J�
�Z�!����zC;5$/������~4�}��?�/KCK/��;_�u𔑬0��U����5���(�����{F@$u'5������#��86�sGl>��7����qz.X�W5�B�vxH�tA��à�Ya&i_���t�7���5�l6�yÓ�<�v�z�0ӆ���:���ۻ@��P/! @��8L./f�u;��ʂ��Φ)4���������mRfd���:p߭�^;<|�V�b������\��O���������� upʌuf�yVC��[�5
�#J��(ɍW>o���~!�<<�) Y�<���S{ֈ�����W'�2�P�K�w@ɺ������Gk��2..�YJ���Dj(�>!aw3P�&��^�.#L_Зڜ	"�����GrS�O,�D���H�J���x��-7��#�;7==�S����P���uC:��=Bxt.�%qɽRD@�{VzG�3���n�U�����0���?;���ǘ��PĴ�;�k�{"��_�=�P�걨,��<e�B��H*p�#��0�&7ϧ''c|���k)����И�w�����閉��-��H(ѝ��j�*O�9�l���sC}��Y>ŝ��2�P� ��Eo�X��,�w�Ar\	Ǩ��n�P��n�����#�{'�q�i
x�"�kw���Po9Ц�;w�p�C�h3�(��}����ZL۽="p��>�u��ֹt�Q���o�[X���=6�]���X�[vYC�usL��L#Ξ���<I�;A<�<�Ȋ��A.-�K�C���L��Ծ/r�1���lz_�����ϟ���>T��K�7z��qH|����"ןZ��JJ��U ��JHg��}V6�����֩{�S@m����{[�l�!�lP��PQ1sV�ꈀg�z��gB��Tb�a݈�n�����Qc��S(f��8���RH� ��%��G�zL4� ��篁� �J�<�;���좦�ݷ���]�Aev)�CC����</�����W���'''9(V����O,U�ʝ�"�W�ܖ((�Ѹ�:=gaa�?��:6��sZ�zX1ݝ�{��o����Q�YQ� ����Y�4�B-@�.���rP��OF��L�E{2��+�	B:�. ����2��6f��L��z=�>I��,I�~��=8a #�ũ,�}fu��Qir񰶾��ݻ����+.w�?��o���:��G��Ȉo'�.�a�d�%�T� ��T�`kKg\�+^����)E���ghXL�g"mȐhHw��7o����w��[��LMɖ�>${'���U"*�x�����K��9<:��)���m;+���(��)i��p�����(��M�f�>ًv�xs���H�!��`f�`F�E��\U��>�--v4obz,���w�I�����Ñc������p���{�(J�c��G���-}C�[\m�Z��f��H-�[I�"�gf�il�>V��uϰ�Bs�33X�RsS�!Ob����gi�N\\��c��b8:���ݔ=����͹5�6O-�8$���/�cьw/������<�KNa{X�-��8�s%h �Z���E*b�>�b-h�R�W�*�fd+�g�H���n���G���H��������|t��!��5L4�B���dRVT�W�KZ<��a1�4� Ղ��<��@R-��b��(�g�|��</�fo_̯������o�wx���7���Ŝ��}� {���K�ȧP�a�H���A������]02�
��˶�R� ~Ä���9.���F�d<�q�) ~�;�DJ>"t��lc�G�Y�o������1�@�
������?I�T		������{����mݷZi������f���	��p��
!!!�z(Ԇ�~~��o��G8J��4����q���D�%<����L*f�r�8������&�����v�5��iL�y��W�)�F^b@|����z�7HMҩ��W�Z;<�j�`�%~s]��{���Jc������.��c4BG�ȿE�k_*Xw�J2.6Is|�k�؋<�3-��̎.�]ў��v�����.>����ohBh�k�[Y�<%FtE��3��{�CJg��Ԃ���o��ǫ�+�؟�y�AtW �F����M|^ޙ��SS7��#��Ǿ��� v#3����Kߖ#���2��^&�%����^�2k�>!��`r�Y2����i�������[U$92X%�\�j
ME@���80�kWHX��W&��kݽ�¼��_ī�d��Ū��B"Y$Ϊ���d8��AE?�'�X��"�,�~��goo�4�#��),	�����M��}��<o��Ѕ�/i_��YL�����.3iQ��z6xǨ���?��-5ukx�d�XNN��'Hp>=l�ސvp �,xm���>(��e��f��d8�PYu���c�6�x�:R��y7}��±E ���������נ�5k�ڋ�ZE�p�=���Q�,��8���p���1U�YJ͌�L����w3�PbW�����k��«ޕ�\�h&����O�&�K����0b/t��o�QeiCYƮr��j��;��d���}�&��u��7�^�iq�o���,�)���_N������g�E_��W�b�$�I��ژ��m���&S��|I�uX��l���� \YˬB���]r�!7<�D��ǊL��(T�~��[��Ɛ�ɵ��(�&���S�J�nn����o��>�{�:-���U~{�ny�^������m�XTT���/��Sy4:���Ξi*�=,�^<�:/���'�H�������6��ϮAv;��?�0ߨ�.go�yV4V�|%��x����}q1��-A��@����bח��ß��,h�J����뇷���kƏ�a8@��2H~�(U蓪[�-0�=�H��!�������Œj�-52��Q�`��[��Xpz��F��v�6Y�
�6�ф��,[O�g���i��B%^����-�N��wBd����X��y�<�wW�� {V��nDV麘m�q�5nM�Ϧ-Z�$����s�<⑨V�6O�%9jr&P�&ED�7.�VWq�"��G�gml�@m���ojo����b�:�FB����ԁ>{��'����o�*�(m�K4!�q���d�+ό��>�7�~��9f�^Y�P�?g1`�Xg�% ���߲5TL�-s�9�E*��rx�Z�LTJ��7���%:ߙ��%J�}y�`q��u�kSS2&�|?�l������
J�ͽӥ��5�z
`���`�:6>5, Zξ<���PN"��(�g��Y╹6ä�C����&P�\�&�,�'&&-��#3;�
�G�rF8^_�O�V����^��=�X֥k�dC5|@5��g�EPU`�~�p����6�~���D��m-����F����j	/�DK�Y�kd�l��QV�gy��T�*w����Y�~-g��Li'(�E��U�Ը6<�ss���������U�w�
/dM٫�5�M+�/�?z�.�t������3j �]E����^�N[���d���!��\�.������&�+22��a�V��"־o��'>�a��D�<`M���cA�&?�I�-���jH�Iy��A1��0��,)��mSH��J�/���<b��Ukb�(<���~��̷�w�xw���`9:l���1hWFmʡs:05���׵e6tlll�&R�D ��[�H�Dr���V���F�����ӄ�.���Mhg��PR��?L�e#���Pj����{�j�e-�b��V�������3��1��'�
9���=���\����A��[PDw�4�$���ݼu~��i��my>��͙1�~),/SoH�.h���tf��� S�
��s���b�(יl4��$%T�Ы9�Ǹ�@���G�x`fַ�C:��Wmk�½4����S��|�K��/g������!�X6s����L�
C���Iy��naӢu�	���p����ŰB�~n��PH��dU�g�5&[����?�2jy����6V� �_S�9�&��&Jt�v��Hb���C�f����V�C�>j����p��"��/҅sD�޻kY'�19LH)_�}������bJ;\�]"g���-��j�]���!KYYni���]d*n���c�(�w�����-˿}���nm��K��E ���Rq�y���}j*=��{}P��] ����Ĳ��û�s<6Nf����[��E��-Ȟ�e����R&�H�%�}���>̀ ���c�N�޻���[Yy�ߦF"�@$���1^Q���wf{l��zy�Z�	�N��2cj�~�%�r��Llu..~Cذa��=@�:CE�M���ٸuJ���[y�!�`��+�|^NN����aY��Þ�cçD-�V��w�� �}(렙@Y����Z�ų����u�v"��u��->�gu���
dj?�ɉ����r��9ƞ���~���[T$���zà�(��S_��tsy�n�7D��q����o9�����T�>����Pr@���X1ȆN�E��0���M�PyJ���_��p������/�ܭ�P����IrR/c;��09$c*�&��w���)�Ԗ�('%>ж������{�������\��:F��[�r7�$�P��o�/���O��9 W\̝2�y�U�Q;�x�j�nP:J�IH,�`��/T=^�wp��uμJt�D��
�������{<R-$j��*�*����,�*b��N�B�������HYh3z ֐��)�ƵϤ h5�����A��Ik�Q����e0�3���(�""8$�I���1�����I���O&������s��힟/="
���}�����d��'��&��2�3G�f�0����s;�ԉ�"
2�4�ƀ���Tt�K0����1S�1qҍ�=��r�Łv)���O>����&��66V���C�e�nP7gޕb^�	�'���J���IDF�fs83ֿ�x�&�7d�W���~3Y᧞�=��n�('}S�f�h�	7<�Ƭۈ��H�P�gx�c�Y}_�j֜]�(����cA2"pp}%��͔12����
ä���d{q����HT"]*���[N���w@r����1st���[���NJ��㶵���w�(�O�A�:?��U6N� ��|Tc�S zǈ�|�J�!Y�zidA�[9����.�:��i����C���!a� ��b���^���=k�nQ{������J�s
Yḵ����8Vm93�P��{���"�s�wN]���)I����������6I�x������*�r)���&���ܜQ�����ty�j�`m�#����9��/}��NO�+�]��/q��7,/��v!�v?��Ս�%���vpP�����\@�x/
�Q쳖�z��*�Ez�* ��YX�F�d�ۀg�E#-,0<,�030w����a�,!�}\I�4ᵶz�Ū�`�Vʉ������bh$�О�
�_Y�42������+�q&�i(����_Mv�9(�F����mU��}Ͱ���ۃ�G���V(m�ti��� P��!h\�:IojlD:]0~!E���:n�N�a�����I������8�z�A���>��#�������c�%ķ�����_�m]�}����p�;!�f�#S�u`:f	�����$�Ps'������د��F~b�a|�-��Qm5[j)/�p㖿�Hc4`Y3�1���F�iio6d�~����M!��l�-��s�}9���c3́%Aei�Q������5Z�a�ݯ�㥩*���S��SSߪB���24�G�r_�[jk���I�dƠ��"2��1���{���n�'��|�Y�MSG��jo==6@J���Sc�M��7f:���MG)�B�v��a�Z�K���׺�z�q)X�`�`�1�-[6��o���=�Z�+ s3Z\�rKOO�_2eF_Ǿ�;��G���O�.�"��Ǌ�a�,�s���*[ ;��j���|��4uv���D���4�q01$�O��xđ0+oi�r�%�|vky�b�����sZ�:����}����KY^lH|�6��&&��`�FCTl,��g�����YC���zC]�$�y�Q���l�����-��H�u���`U�����+�����o�4"��6@�������k@��$M�}.�����]=�z���𜵵G�=�R��2��Q��B��[ e_XJ�bAcctoo5`qqE璌�"�����G�u�<O����HP��d�.���g�mlp�rßqS.�_qy��p��l��ݻw��-
u�k蘍��oP����۰�����L���I���F��� ��1������CX9�~�xP6�B9tSJ��i��rI&�l�6Ǣ��>�4>��O@MQ�AsRs�u���8�8�s3O�
�{�=������Z����w�� [�ҴGɮb���t8��_�<���C�����~�nm�e���z���Xq��@[�A�'50@4`ř��ϳ}���%���C����v�]�2,H�mo;y5r�남��9�ԝ��sQ��iV��'#�R�"�*����.��X��i-�AFjI?�z�o�ߙ����
l�J
w���5c�e��>�7��n B�Ʋ*Ԑ��U�{�J��/��{����BB��Ռl�%i�*�)zn���}�
�~]���ORj��(՜.Ob�L��}�^�]JpggHRJ�.��5�B;*���6"��p���9������U^���S�r��(��	4�"I��k�q�!q����bs~Y����)�B�6�xꀥ��C�u}`Q�'�m�0;�-� 8��]&�[�S��P�x�nR�{��:�� d�Ø���)n�ܸrK�0�o���ss�6s����;�s����C��h�W��0Y�QbvvQ��ႉ��k)iiHd���=�&}_?AB,;�"��8|�l�[ظ|��J D���|������-���9#uG��ffO^h5�;(
5��^�W�����Ĥ�P�N�k۳j5Rp���z?����;�� �6P.�s���5�-��8e�}����xJ?�ǁB��#�6�g\�q�!"b?+ ������S��x@����%/}n�M}a�9<��9���`�6���~X"3�iJ<�|D���������I��	K���읚𑍎���j�sߵ8�]]�Rɭ���X�]\\|���a ���$�넪��S��z��/(�jY��|��C�`s�����&؛E�����=A�D�*��}�"���ރf�v��%�:|����Q��QQ>��0 %��t��Hw�,��! )Hwww����,�%%�������+ҝ>s��s~���⸰3s�ꚙ���*��8�&�y��{�y��s\\O�6�������1����j�����e����0�x}�����*I�۞uNd�ሇ�w��W]�[���E�|�+Ra��G�iL����-�.S�1���:��8��+��:��������K�3����"/���+��}���^qo�~|��X�}NsɝڵYՈMz�mN�K�m�����tW�B���@H�c%��"n߾psY�qޙ�$GF��C���`��]n�wv���7@��
��Z�7jǿ�Dx���ׯoQO�-��[��� �R
�����1�p'L����ZZX��O/��r��5= �J|!�7�팋��+��_�� >~=�K�K]O�ymȞ�Z=��E~I��e���Q�7��ygg�s�7�888�E�q��u��}9��_��dC@D��*-M�<��0� X&�zC��jO�e�80��i2�����H�߮�#Uw)2�{b91V�c	��^ ՟rQ��*������Η_HT�Z�6�;��ݝӼo�;�v����o^w����PQ9a����(
�}wP1�T&�
+*j9n:,2� �RsfR|�
�W�O~��3鼕<�`i���`���KY���Ip����c��������Ze�����I/�V�z��WdB<�,�6��(̛�b�w
�����cE�	��1AЇ����:le�p�����TRq����F��跉ec�;�F�1��������o�b���Љ��m�f�D���Y�����ֹA��(����yN�|�53q�e>�͈�s:��iЋ�x�'������	WW������A���G�D�L`#Ƹ�(t�@x��S"�uV�+�����1��H��j�&�@F)Ϟ]��*�B�I�%;O=�H� �c�H�Nc3�|?x#>�75����	+�
�d!|�ǂ�����?���;R��r�E����,��g9x�hV~��002����5R�lU���2�C������� �C�:��ŷ�[�t��I�С"�\n>�`d����@Nl\��~=0��������70z���	�ۓڕ�/���mm��{Pcٿ�����&��\Rbj������6��G�b�� X;����m^dވ�y�ų%Z��cu#�d��x��v�M��������^���m�s���d�kJH��3Ux&��,{�~�=�����rdك�痡�@[�T@ۛ�.;j��9������趋}@��q���WH���ncj���t���"��vh-+k���-e*#��а�����?�XY|
�h�t~�� 
�"�����l�b1��"Ɨ6���f��m��%�\�U�ŵ�4HY��������u�5�t6a+��o�j��b�;����ȝB�X����'< C^��N�§������p�^����w������W��7	
B�t�<��w�~��_G����̜ǭrh.d������$b�#(�:��ũ�3������!�����:T�(rپzl�����؈T�U�MF���`GEv�����冷iS�s>z<ݥ���v�×�6����=Iu��do��K����h��P��y���hu�`0o*�kn"Z��Ǚ/���	������'ѹ�|v�wT[,�*%���5�"� ry
��>�(3 '&2m]]��p�vMLp�D6n}�R��k+zя=��r��xe"?-5u7`�����mͣE4j-����6�ijn��E�^	�U(��96�NL.`.Ҹs*!�c>ξ_�@H�-ͿΥ�rs������%555�D���k�{���]w�=�i��B�0FX�>D���f��hb�ͅzyLR�l�=���Y��p�'ė���Η�|�Cߵ��>�����Ed�ںF���Y�{Δ�,3�)����#�wAM����Z�Р���^��ii�z��������mA�I�I?���}��n�~F;�8�ba!�/���{�ϯ��x��v_�+�nb9��GD/�w�,~i��X;8(�N�hTUW{�����&�x�����|YȽ�w~?AP�%r�rE����б%�"1�ھ|���] *�1kZgD���~,OE�0�}�l��C�g����~V���=���&��N��hK�LhK�5�<��.u:��KD�HS��)�"��oW]�����4;�dI�|�R7U���z�֔�:$��dm���ǏX+��f�<��~���ܒ�e@ 9y���
 C�X�������_����� 4�y��dNd���u����{�۔���s?�-�A�����Ò��yv���������v���cz��O��fr���f����^K��k���)��2������$���p�Õ��4�IW^���W�	&	��7��g6$��­���]'��m*3${���//C斗�Bca�����>����Eo�l�P�|q�ւ5���:J, D�R��w]�u����ggPg�чJm��������8���)�ôFl$$��ղ�ˡ�Q"uMM�elXᅅ,�ĉ��}+}�C-�HA�qS��qHk���Ņev�� Y�3�bVNL��⼕Y�3+|�?��~52ӫȷ�{k�L��lJ���8Ą������_=I�x����0a[��.U�{3������\���-����PfH�H@SK���f|O�Fsy�h�FUMG��v�(������w2�|Y�!}�O<=�
�KQ����@꣓f�&"&~jn��Ǝ+MEU��w�d�$edꌴ��avT��@g��߀o(*%�|y 2F'FKCV������IDH�Ch�+�=����𹶨g�b���.Y��3��}��q�?M��|�u[�y>Ҋ����N��<�(���	����e�������,@4�
X��	
�:���ǣ"g�[������K�����XU�0Hs�'����x�,oim=�w۬s!�����'�/?� ���_��.��1��%�y�%)yiy_�e��aY5'������a+��:w�Wll,do�9Ҳbt�>�R� /���G�����/��L��$JJ˼���A�gV׮-�=��-��^�.����~�&�� k��K����7�r2q',���[F�'8&~�_V��[^�C�dk �|���e�Lg1���;�Gw)��v��"��9���==#��nWyHп�I��f?6����H*����)_&�������#��O��?AY�:���+~֘�vD�݊��O(�����)CCFĦ�'q�	�ܻ뉰\M�9o}����.�������)I��x\�n���];�(j#����U�R����Q,狭d���ֳ�������s�C���;��v˥F��8Cq���	:���DuWv��;ᨯM*0o/C⡧w��?��Ȅ�T]�U�	l�z��%��'���\\\���%UkDe�{��&�0ɩm @�#�ĩ�<JK>궎��i���S_��s���S�hδ��1�F��2+���dm��PVc�t�l^>���<	��C�È՛j����ن?*�����{p�-�9=�Gؚ�v��e��++lm��G"�YUĞ�Ƈ�6?�
u=:$a��
#�ĭV8�B�ry�C)$0�龮���`�����V;k}�o̪�����w9�R������lh�i 2i�ث{��*F�/.f��� S�P�
�w�y�V��b�[��������H4���.�y�H/$�3}+���k�30].����Ε�����נ]����{����z�8X����l`���tTҜ���3�b����%?���@��f)Xb����? �#���yh֪s����$��=э�[��~�`	dO����q���'�d1���Q"�=/�~����d�a���uT>�1��	 �9������:�Ur��;qp|l��	��--�^�f#�����[�hSp!˄�7�'�.|��hl:"X��fb��P���Z��&Gk����(�� Sf���
��-���g��d�!!1��1!~�����R��u�W��֞��1S�얠�t�M���d��M�Y�p$��Ry�#�"��j6�P;wF;"N�Q�&���`��.楫&�遊�m�#'#�9IB��fǖ��[��#�/!��QmR�=_�ɕ8<��R2��M%�Ð�lEmdf��n�9��#� �%L�/�!�ZŠ�7���e���$�Q��a��ddf�%  �������{����=_�I���I�x/�����8��3o�æL,6����+���
1YY��v��<y�����.��u�g�=v/���KXh('�ꪛ�fm������W{�#�mZ��阙'N ^�^0���o+�>A�p�q�/�62�Xh���WM��R;��:ڶ�Y�n����NM��@����Tѭג�,�~��Ti�}!z�`p}{-���9Osi��Xz�?Yii�{wщ��0S>�&5�D�ļ�"��?P�W�8ݥV�r�g=?<<4>��ZBp"�G�B(`d� $q�_9�@|z�I�v]�E�ynz�I����؜���ٜ�+��k�}
�!���Ǚ�0/0����m��6����`%���qP� #�B���4��� �0�<�	Bb�=�©��o���Q�0-�4�����>��7��M�ŉ/;����1���mϬ ��WI���o2>�q�K��ɪD[�o��������d}����݌�JLL,i�@���'޵}�#�Y�������������zK|覫�����Eж��d'|%���)&\���dA�U�'�83a	;r5��Iʇ��Ȑ��1���lП*��rH�橵+�xP�bc���-��ٯ_�y����wŷ���>7�61<���h=�J�������� �dȨ�ػ�3���?� �>��Y�~�CL/�a�$N�|�i7V���GE��SS�����#�ohj�C��Q2cA��J\�Ѯ��']Y���w"��L��eX��=*E����/��*%��͝�����˗���|����-,��#����^1�mE�>�"��@|Q{h���#@�>h���.)-+�7��|����0o4bO�y__��49S�t�&(����
2'������QT}�� G�_���eI�������J��o��۫���.1>\nmͰ��mE;���;=]���!}�)�1{vХ2�k��~���pC�����O�:�}_On��V�'H@Q�jAs��9t��B��Ԉ�O���_���������"��>^��a��_����e��z�
oi�v�R�rM�VM0��*�kYOwoo��svZ��:����9A����#g��r�VV�,�?�Rc�Gs&(��`T��?��J�Лiq��tO��}�����Vi�y͆m��-t��Z��PR2v�z^��k?{F|��DDB� N���+�� =}���7�,����o�Y��Mo�R�~_��_׻�~��8�`�!/�z����OS���2��<5�3��8��z�$�ܰR��9{i��Ü�2�a�gK����d�6��Z�Q�Q�UGp+�#$Kޞ�.�e�Ff!Q�zr�A�����j����1/��S��ՕQ+_&fv��NXNe�8��$u����#�Y�P5���^����>�<Ɂ.n4sQ�,1�rRXC��:�cbrA���^�Cvp`��;9_&��9P�}��;y�Ԅ/���,�#5�w?8<���p����%���~]ږ�_?�h�IB�`b��e��i5=�'�
O��k6rݫ��翺��5ƌ�49?�｜<��^$"���$�Ǐ_]�Al~w��Z��-B�1|� G>��>�&\����^�'�6h������Z_�*o�/#�7�����0VU�D ��O���,��S|d�ӗ�-��w�EA �PRQy���l���+���Z�ww=�[%2�G`��@���$�#�͆��{�1f�jv����σ� f���l��	��8h~�������W���5`他B��I��O��i�����!����=��L���(��v�Ŕ�/ŃMe�_�.	�JW_����:.ٔ�
�wk���׊�S�JEEȇ���u�u?��ؑ��.�{�K�/��"�&!'�;z�X:e9�j�����
��+<�IAaa�*������i11�*I�a/��-�ϭ��;��t�ﭜ���t��j�s*WCg��*C��x��X���Fv�����XV�16��[o�_]�4��Q���Ȓ:����_o�q���-�utxx�EL�y��[ޡ��۶���ᘥ�/ֽnv���P�w����5������^��2w:��H�4����(zt��A*#����iq�>yW��n���%���/!�����P��v��3_���jW�S�|k{RGmʷ���OA�tR���d�UU�� O�Y��_�nRi�?$b��ikߌ'��g�V��辽L��MD�O��N��qS9����U�[���k�f�پi.��y��<3�Wq&O��\ڷBo�UL���[<8B'��s��-Б#o��X<̶n�t;˻����FG
0z*��k���X8ן�����0a���Ne�iAp���i�g�k�uz?�\�D����z���Ȓ;s�X~������h)������[N7�	!�2�3��ٔG��u�K��+5��۴_"�����|q��'Yn#cq��h���9�&�<��۶,�r�_��`Z�c��e}��~oo{�o]c�g��Ǥ�'�09�-��_�XA����;��q�����C�����.C������#�i�_�n$§h	q�x��N�Y�C��ε�U
�5�-&�C��o%fd��+���95t�,���C��NEm/�>���}��ݺӆㇶ	�`Fj�ɺ��8�Z;Z:|캖�,��܁U���T�Z:�K�1tOmO�GJ�^ּ�v�6ō,��5:\�g7�;�T�/�e�++��]`t)*SssV�k��X�}���Ԅ;��	�4�T^^^Ō���II^�*��-c��"@��ו�M��,0d�3���42d)T��vy��F��)?��S.8���8�v�iX
�|u�m�ǚ�ƭ��C�*�-πmQ���p=�u���}��N�}���l�X�߿��<��yI���Q`������pcjB\�㭠�B�I�+�Ծ(���ۆ�&����ɐ�}�'㵡Q�����SW�%/��;����umE��m��^8�8Lͅ��(q�mk����N�.��4���ɉ���Ӗ��[�LII�۷�i
�x�^�gO�L�M�;���7]$�w{%�GPay�v�S���F���I02��@O�.�X�Q�#E�[m���r��\OuUA�����Ɗ��������4ˁ�U*/���bk=�]�sPz6��io/Q�:���R����8;�#"Y�_�6T'W�E�?$Ŷzpr4��p��ZTzv����un��G�v�򜁞!$�$�"st����3�4)b�#��XI>��&�����=�dqi���������P�{(Ԉ���Ü�5%fR��~��$Ԧڋ���{,$9�s⯢'7V��aK�_ZKfƟ�9ã,LpP�Z��\��Ɯ����&/ػ����B��OW��n�UVpwK�&�a�ݽ{7�R��%Tij�ǃL��1�Lx��+MIONL�&��|I�-�v^n۾�:��Q,'z:ha��2K�S_(�sm�%]4b��Ҵ�����\�@�s!us3�������J�&� ��ޖBG{K9k}��VAߊ��x2�8���>�S��!1��XS>'�}+W���\;�
ޏm5d�{���(z�1�9� 
���@�<gG��e�9��L�8�%��$��#�k5ߓ+6�aJ�[:<���		z�& +Re�� {�W虘4H�X:9��L�{��RUe�y��-�Ք�����\��d�,��l6wv�����H8f'���wp꒻@��Pe��@YdH��)M����|�(��J<
���(�0�ş���*LJV��jr�uVzw L[��o���
(�Qm�m⢃���l�]�e�ӝ(��n>p<4�ʻ���N��C8r}j�>�Aqn���a��g�՛�@�� ���%w���pVn����1������n利�?M���+�sU�PF�9�df�M)4��S�J���ȽŴ%6d� >�y���y�V#C8�.�%`�ݥ�&vf��ꠧ�LFkA;q��������MϠ1�n����3l+�\��-!yj�cx`�ɒt$�����DCs�� ������
ۼ�VRߊ`�Vn~�J)�=��z �''|��P��'�zm.���އ�'r	�$�k��/Eғ�i��|��Ԛ5@M�s��Y�i��=[lZ����(�_���㝜�N���i�Q��^c9�8�>X�9Ig�j�uQ4yP�$
j�ZX������z�$�yz��p<�o7�X�����+��kE����Bs��S����\+o��#�Ѕ������gdİ������軷� G$��Vu��x���d3���4�6%&����B��oL��$B��!��R�:az� L`�l�q�L�8��gr|�a"����B�	}����or���Ń�^��E%Q>UJ�2gء�]+9�C�����!���OdI��^��������B�q�x~�S�����]g���9W��W�Č3 vAdr�9�~�(CX2 ��[�x��9��0_`�:�J(mT�Alָ���xr?�gkce�)W���Q���n��Ut��ɟ-���$���p�Z�_C�w ~-8{���ϥ8W��7�(�Zh]�5h��s��u�6L�����ʍo�6���^QR�ԭ�����W�r��L���$ʏ)*")�|���911T:�v��n>mǈ!AO�1`��oN������H$^ٯ�DLJJʝ��L����X9�`*���-.�[�q���a��`�m��i�
�c�?�*����/��D����6�ʰ���qF]]��#�W�|t$�oФؘw�Vr�HijI���v�{K��O9h�����6�&K�k��o_�npa�d�I4��j.���y�)�AoR]�Ph�݃^BيY�g�������=�S^.���&.���(S��{�u�l�w޵�E}z�F��ٲ�k�N텳�����Z�w7��,�7��$Y\$nT%�3�����	rG��wg:ն�����ǹ���5^R�2`T���ٿ˹�Gq�.\d�W/������,��Y'	����(�����|��f#���($�+z��I'���=c��|����s0��	nE����1�C� t��ȓ����r%�@���E��qKܜLK\���C�y**a�����U��/nmz�>,�Cz���k���Y[_�w�x� ����15qJ���5 ]7���O��.�껺bT)B��Nl.Ϻ�E�HYY�t(���;/Vk�c]�K�3�.��:��M�[,(�?��p���[h�9�HT)22���e``�r݆��?��+>wp� z}X����iq�^}ش��h^� �×� )�j��s���X�X���"�]74r����m�T�=X"���ź�O�����m�g�������C,x�k�\��$����Ms�h�ۂ���t��ܰ�[c�PL9<�65?ˌpL��b��o�	#╿�ʹ�a��E?;��)�,;Ҟ����2 `���#t	6�XUB�r�|���e�v�h���JQ���Z/��+��
A2J�����,�{� A�!_k�աuw����T�C�_b**�^I�$�����m��a��E}�D��ׇ�R��8P��pvu���C�5`�4P"y�'�+��A2�?<%�iI����Y��Q'h^�7�<��gfEX����C8׽�2}>ޡ��ʑj�Z'�ӑ�]��v!
m��f��^V9�����F��M_��{/���� R�lRbE0�\���R��^$ҵy��N��67���罽��L
��ϻ������뻏�b��W��B��N�sv>�z��-�5��vQ��ܹz�C�׮��"黦&�)wz��%��Y�@�)렐��8�
�>A�LgX�$~���~�s�}ޤ�ö�~���/o��U�s�r����T�#֒�l�JTc�	�����'�*��k�J|.����G����Ax~I�n�m�׽��u���OU��@���3���t��u]�G�<ԝu�Ŗ�{�;b�p)ǭ���ۢ�Ti:3���� �����]r��+���xxT�C�s4�Ss$�K(�8A�ڳgĜ3{0T��S�v���))�KF����N;<In/� �9h�(~��ߠ%FdA�\'GM(g��|/0��	�Y�5�7�f����n�����Y�)eQ�.����+ƪ7\�ZZpl��We�a�)���� ri��|!���h���/�����T&y�v�z!�O���&ݟ`������32�U_�Sg�;�cc�X�I��x���P��E�����mY��$������3*�5���`��J<��T�W�� G�Ǳ�h�_�n;!ȌYҍ���tTJ���D׎t�UNn4��ކ߭��
���ӹ�y��;������o�h����ᑥ����P�B*;�(�����n\o%֡ #|V`��t�=rӗw�9�i�V$8�yT'�YJ>�יN3
��&���\z���؍���\�5��X�Y���V��(�܈���̥%�q�">6iO�EjkZxE�}�q�L��P�ߢC�5M ��L���-s�	��<M��4cJ���˧�T�=?=�ssݵW�n�ߜ���E��n�<���[�k0��a���^�4+P\��jhz�Ʊ)��R5vG��PϽ�s|T��[�����vy�Q�Y����;�+~�)Cs&��7�g?/q���N�O6l�<�̚�3hmmc�s`�Ά���X� �L�S�G&œ��o�ί}Y��I.������\p��"����ܦ�
.�vh2��`��=�$�D��}͠rV��B���� G�HD�ƞl^�7��
Z���������@�v��'u_6~If���u�M���Ǔ0�=�dk�?AFGd��qm��������"�ڥ�5r ��ÛLهa�**$d�C��V4,_>�]��p�=��-��lNY(+�-	�֝���6f|6e�����;G�|�{��٧���?�~�ntӷH���ō�l��O�,���)u���M&�%ni��$#$ͳ�b*O�[9^����v3!�B�:~�g^d0B�~���ntX'p%�MJֹ��W$z�$�w.��l���$��� ��@��I�Xr��u�L����i�����X櫻D��.�\�Y<`�Bt������.v/����Y
w+�J�}��jK��X��������hv��E}%��2�|*l���Y�1��ϯ]nj���b�u!�ܑ�ud����:1L�����.w[@ظQ��&��#E6���������3z���=� %�i3C�%f�x\n���b n?�/s0�����~��#k�C�+͋Py ��M�X5ĳt)�/����.��g,y�h�5�/�TV����9J�~-���J%
o`�ja�H��J��2��%߷�ɒ���>��o�����*ྥ�s7���)���c?��h)�,ʺ),1�f�3i@NS���o��-�/n��*���}dJ�F&ff�P�&���F��4���z]�Xk������g����v�q�l��߿k��;�%�^�q��CvlR���B��O��*&���UZ+����ţ��Q�j�2��2�u���@�3����Vp��Yy�"�`��}�]���)V7�ѻx��\�]����7�Z��*�P�X{x�0��]�I�W�B��W��-��CMY
(�_��茸W�a��� �0��ܵqȒ���m(�v���F���d��<^9	��9��Q�8�v���RҤ�wM����b�����㋶�Q���;�7�}
���=Ʋ��y�j��������4�A���{` ��\�����x4p���hϖ�'u�V�0--�,��»öךLƹ`�"�����y�:]QP~�V�P����p�l�X��l�a�=�*y�C��>um��Ζ�C7.��m)��7
T�N8�cI�9�n�_i@�!s����\�k��m.
��Xx2�@�k�I��U�O+�ٽ��X�cmӕ��5��o}s�og��Fw����R�C��#u��*�[�������C�]���B�#��֓�%��RN�^Z��я���Ε��x��qNw����>��UW�|0�=)�/xc�ơZ���ܵ�b6��\'h3��I�k�!$�����V^��~��
c�������j��Q>��M�И����cn"���a�Rd��✌B��
��Up�jR}��E%��Q%��ݠY���h򾿌霬R��p��}
e�0
����Q�L���%(���^{�_(�$ƈO���r���7 �g��`g� ���;��l��	�z���><�߂-Mm�D�և�NIyyħOr�s_)<��qQ>~��C��s��K��Ӌ���˼���au\w�$��� D�vs���8g����b{�D�!x߁�z��q�u���sr|>c�|���0�2 ��ԕ3V��:�ȿ������D�,�I+�n��Y��q�bہ�9>�;w�|_�7}��J�4����Uw	���(������R)JQ&_ �K�D�&ZN������2��h�P|\���	����g�2�� �����|
��_a1�͋�9�cu~���Ô���tR�=� �ߺ#�2��;҂2R���ߧ�V���f<�r>q� ���"� O��ռ=���lg	c�u^e���x��q����K�(E��XAPh�mw��o^G���.��\ܫw�fܳ�1x��G���������lpmN�"ҡ��U{af�������/��4�*^��q��K� _����5/�w@� ���`E` ���f���z �/3 -��4RB�����'論��7����v�Ɗi0f�uD|�{#����L�R��S����~on��x����2''����3�X�"'�dnb�=Z�u���\Hjh���ၗP!%%%�u�8���<����rU�4Zn�y�2WT�������P�����1'�Bnw��U�/�P��]���wA��|����:K�w��YYo ��6��/��mKY3.x

�\F�w���>��K����v�s+$m6�WR�l�A����ÈF����EP�(g�ZSdʷ��,~��3Ǧ'��F\����B@�?��<� HJ��F�돕]R8����&RL��Ǐ��4���USP�M���� �
=���F(&%����Ħo]þ�g�==��T�%��G{J�O͇>5�/ېZy:�0��[�n�ZZE���6qxH���r>�����"�g�6$��ʒ#+.�Ύ.p�>"��
Q���N��xk�}�f|;��(�d�����f|m�[`�3�?��%�GքMu~{�  
P�'��Ts�7.Ed���{�#�hZ��L�X�Dd>P)�E(`��#�H�gc��|���)��3�_��	��Wt�Zt�q\�I�bt�m����W�57���)l�U*�ck���d�!�zR["(�?���t��Y���7"9���~10��A���6�ε�ol���u��.Ri��+��_ �r����E�6�K⦣��ra�z����:*�wӍ�	Pŏ����:��;g�{����qH�t��\k,�_��q��a����'C�I�ꔷ�����ɖ�����#���s59I�x�r���c&��c�ǒa�'����L��	�vG�5w	f���[�X��?���@��X	�c�'�N���5�c_һ�̿]P�:��Ԅ�(�`o�u���1���A�M���d�˰ 
C�6egu�1		Hbے�vd®��� m�mw�y��1��JA��ً|��U��;���g��je+7���Fʙ�)�9>���(�u
egWW������?<�o4��t`�3Ԫ
Ş	�m�G>������z����B���ҭ<�a:��c�{0l���'V,rG>�黑w��0Nɿ�V����sJ[�Pr˻�6ƌt+�R�Ԅ����Bw7}o�e�z��[`R �m���M��e{�0	#x.r�^���*�O�O�d60���XPrz�"��J��X?��j���¨�������܂��0��@�֯.�`�P��ɚ�Yɖ˺���� z�,���#̑��Y�4��թQ��T�E��Ǐ?|ot�\�^Y)���U�շ~��8v�/��*�?��*EH��_�SJ����p.\�� W����z�5�N���fM�B��TOȅy�����*^{X�0�*>�+\!w4 )u�.���2d�J��IkY��8]��[��a����9������:_"+V�Z��/��O^/~���F&&�?���S�rk�*��L���VMa2 ���l���W���{�Ϻ|:B�c� ��F��EG��܈ݭ��?Fڋ�RC\l������3[2�OL|4u`1<�uj�e�/N��w(�E��Ӧ<�q��`Gw����͔�3�]r�I-���F���-�j�E:�IH��7.�82E]��_��V�"��*��]�9��qǞ�C�}@�tTY��Wj��qQ��U8�7�j	�a*!OW cj��<����|�aƗyi5�B���SU*/vBԏca������� 2lԄs��P������\��"}��H�--�m��J�;g%�d&��z���RV<[8NB�4f�q3VE���fd>"�X�YoLL���]��,���g��ơ��y?O��<�v�8���⨾��=����BO{�z����b9+V�fi�>7���cô6�-�H9)��(��ˮu��	6BOO,������7��`f�?ִ2�\�R8�`�a%�S����z��A��>'�M��.�G@?\F�d����)=�r�Ț�GJZ���M�|��cJ�}����ɐ#ױ��w�\�7���Y�sؤ(A p�ж�x�ח������S�eu�+}��p��LǊ�u�=�%�J\1�"���e�"wp����@<���נMbݳ���+�Ş$"��u����59U��"K�hm.�u|���?�yp����Oѿ�ĝs�#�M��䶅"��5kkS>q>�A��z�=v�Q7TǦэC�!��PC������i����:�60S��Hg���&7
QVd��u�M?����\#*]�������e��G�ܨ�y�qF�V8�W"�J2�����m<ϙ�A������P�xlL���nN��ߝ���KYQB��`0�ϕ�j�Rh�3̝Dh��O�GSc�T�im?�8p������S>���"qu�W��KAW������4X����611Ah]?}C������#���q:�$��>H�'�)�l���'�q��o�]b�n��W)V�S�9� ��-�CFo�z<�׿&X�����ǔNb9FFF��v����`Ry��C++YhS�4�xpejSP��P���C�g�����PgD1��i�_�P6��e���8n'��9����A�8���Pצ/�{k�y�^���o_<�]�.�0Ƹ9�����
�S��cɺ<W��C/}��s�ڤ/�`i���hjiM/^b���~������%�.Q6&� $�XrO�/Kz��Ǚ�ȧ�S�pf�{�-q�P!��j���Ȳ"�Z��u�j9�2�q��Gtx��F��ň�Y��k^Vx0���n$Ϲ���0ie��J�����o����7�Dn��r�D~� ��Z�~�!E�"u3j�P؂�$���,��}rl�ϝ���sQRW��I� 3�x��lh
	qwCJp�V�#1@���a�@5���M6����kfƫ�֍��P�k�LQ( ᥽�!'�V2`�T#�Bp1�o�i̥����gBw6e���(=C�;��B{���Y��!!	�|
� M���M���Ǿ��,�8D0ӈ�&���52��(Ħ��O��]MM�V����A��V ��^svI��T>yv)��W�[�Ī��ƣ�9)����]ϔ���KƏ�� O)�>+{/f�mDh�$�YiSh{���>̹�̐$Tt�]mh�0��]��z�֯C�X%bYx?���o[��XRh'Ij�u+��x�aִhv���V���:P
BY��܂"��ɗָGOw��J��w^fx�G��Ϋ���g��vL���d��jYV�Rr����.p⸩逾��x]+���+N���l�s��r�pffF(o����Dي���X��;K��d� ``����K z�j6���U�F�(Hu=����<�"�����DZ�M�Y��<�ҵh���_)=1g���5Xq�L����b��0'�pF��������=h�u���%�ܤ !j��B�sleEJ�a}[���{�Ն7.CG"�; ���i�O�ho`���-�
E~"�	�[�����Z�|80%SSS�Dh����0�r�C{�H�����Z�x�_��'�Gސ����fU��ǀ}J��A��
.?�<b�1���ڇavӿq8��ЦXyZS�*���<oT]]��|2����/9�l���'?55Z��H�7������:f��F�����1�+1Lo��}92���������/�&n�IuF��p�o[���sb[��wޒ
no3qފ��K.�=�_��L��@ܥ�"����Rwr*� F�M���N���͕�C	Tht��9εtv��`ro=���ؘ��x����67g��3%¿{M�F����Ni���#6i��4��]~�˅ʀ��C�Μ� 5�D���Z����]������Y��u4ڎ�<@�ͤ��X��O��m��&& F�6T�̏�,�_���
'K���l FJ�J��m��[����!nD�������`��4(1h�	����S�pm���U�^�"& 1kkg1i�eKK���ץ���%����G�o�_��KDz�t+�T��*T%���Fd��3f$�N���=�G@@�n���=?���4 �&%9�\b��ƚג�����2õ����E�Z�0U�yV���#�
"N)7/��0i��2iiup����g�###�{�ȐǦC���bD@����(m`��bt��Ban�!
ms��bA_�豢(W�T���Utz�x���� ?W���x�~=�W��Y�F�����DT㼏�:��^��8>c<ܿ�a&L 귅r�LH�m(D9�n��F;6?V+�"J�,�ԏ�Ӹ
�fMS���hPRʧ��v"��Ԯ�5���X(��;
���\g/"���!@=l�Tm��,8@�4�~qd�����o�E �)�ou$�4��>-�{r��=���7���K�D$�5L`Rq a��Л��+�[��.X�5+''�kkv�6*�w�	� �x�_�<��}���gƒ ��c���'P�.���������}�ǉ�l'd�	yKƱ7���!;��{dfd��!;�^!N�N:���N�w��/}�����8�D�����㺯��19u����t�OO١���C_�,��ÿ��_�Q7������]�E�&m�F�[��Ũ r�/�ˋ�Z|,9�>gĿ�-�e�4�W�,x>ӟ7��lh|dV��A�m�la�d��7�'�D˃'�Z�dR���><�
$ �8jNDR���gk!�{ 
s��� ��
� �ݖ��6*�&?*��;3�n��.���"���V���B��7�t���T;ǡ�<ΠG���>��^�U��k-Df���w}/HD�'G��u�+���[_::.�t*��XYY�����[������G��,>#G��I|ެ�`vv�)Y�D����,jƴ� <���S���[�B��A*�Ss���;Q�{|q�%������G�\Q=������_�>�Hߩs���V�,��'x��f�3�u��Y��N-��،�y�VV�"�痟��Ӵy(;SUj&ydV��o�z���z��2&���2S� B�W+}��Sj�Nɫ����[}������i :��V�b�9#|�hK�ɢ8�ͭo�g�ҫ҂種�6�?�F�ڱ�]����"�W��l聙�L8�TU p��J])�64�����}5�>ԉR2�WK����߿/�8����L��yt��1�#(II��b97�\; �|���R��ɣ��{8�~�-��c��c	��3j��?�n���zn��4�'�=��<1���Jw:�>���~/��u���F:�%.p�M��X���6y�\7�Y�"��ņɨ�O����Uj���@�%i�]��Ij����LU��z�U������l��i�:�r��Kp�J�L�L���#e��/e������̥����E؏m) ���m2����'�8Z*u�Ļ���s��;i�P;�X���q��^_T��X��:L$iկ]Rvf���1$z�O�v��\~-�:9
���7��(ɱ��T0����w�8T�6��uͣ��˽Ġ&�ET9�����p��wehhg�u�[�wS��?�i�W��&�1�4K^��T��.s����HA�� ����v^:��u���v_Q#q^�`�R5���ܺeZg�]����A�NB��[���-��]��F�Q\�t�?-�lUW����M.��g2���_r�q�-e�ܭ`j/�k@�}�[EE��B?���N'~ GߺN����aݩ��]���ގ��n�rt]��SR�n���Y�?n���Ya�-a<pl�j�<���~� -�=�z�)p�,�<����ܹ�x/_�
�ͰT��~�2ުNZ9,��:]������M��;�t��A�\��Rǋc��3E��f�J)�P�A�?4��+�^j=�rA0k����"��Hw����r��
 �����סR�b��}�ʵ�U�Zet!��6D#b����4�XaY7�� h�[~R5 Ғ�+��gۤC;�_7J�����.�"��Fn��|�j�e��k\?�w� ���݊QW�|f ?[<�#�r��fQ���sM{i�$*К��+��q��)[A(�l�h�e�mp��Ղ�����
��_T	$�N��kԶצ������~�$����w�/����@�R�<�F���o$7ɡ^���#�ݹ��gN��g�+��x��]�h	H�Mh�޽�Bp�ɠm"Z�xԿ�BC ,���)�ٜ��a�*Nq��-��ޭ��>�>�@�D͢��$®���i�8� �2�klk�o���¤�+�.A��g�!��N�{�<M���(4Ӂ�?8Q����5�:0�*�S]�
�ϥۅ�vq{�����9�?-d��S}��r]8��I5 w6>�3q�k���sS��\��V��5�4utD���
9J�Z{x�-��n��k'"L��w�<�&\�U�bc R�M��;>��V�u޶O��t$���81�������*J4�4S��I���z���T��բc"��xi�k�W*���ꛘ�I�G�hX��'�2�=%����Q+uZEϭK�Y� �(~�jZv'����$�~�4Z	H"�jc�g��Tq/����1Q��O����Fv�P��o�X�x$7�,S2���Nς'g��w3�gO��?��wiR�����̧�m�=�e}���ݭ.>�K�}J]P�1e���j��n+R���f@}s�Ñ����b�h�������B^�d�<[鄋Y�x�=++%h���"z#�i����S�kO}�S�+��-2av��ٌ����U��LC���ƀ�|�_~��r#^ͮ~z�Ni/�0G!�>(J'���1��8W&
G5���)��ʱSCb��u��U^[K7�).�Jj��- _{��j���rpx!&e0��^��t�˝����C�����W���^ٖ�Y�2��C��YB�)H���h�n�i�8�����)��� ��{���:I�mq),Q.5X��ؘė893�,-wx�tB�� ��K��-e4dLu"?~XX��s��k~����trA#f��+���@�gty��}��F�ۻ)��Pé)���kJ�{5�zz�WV�	��ou���; ���H0����s��k2;�o�o\�9�QR�v�/1ʱ���d�U�	D	���<�ڵt����S:6
�R'���3���C8����[�uG� K���A,�60����(S+����,(��W�їՂ��N�7L��&�<@�5����g����ʃ�)�d��W���v������~��B~���jI���T@:m�G	<h���9*A�O?�oKY\�� ��b�Φ��� =������)�Ù6I�����wD�@���/H�J�^��as�Ȼ�au*A�6�Hŏ;r�w��e���-�+��:Fg������ϴ�����:�����n���Sf/pwK���du7��8�~E�,�%��Q�WW��Y�l���r�W��6ͽ�,�J%�DA�Q=�L�؉ّ�=�3�7Fr�'��a)�p�tZ�EQ$��굎 �����>햀�*��u���"0K�|05�<en�fG�*E�5q���D��^�;��/_��P�>+���m��u�aa���*`�}�ݿ��ktZ�Ŀ9��Gn�������<�7�(�>6��N�	����㱫o���î���^�*̍Ԁ'��9�窕��Kݜ!G��_�;�7��-"B����<:!+Z�F������z��s}��u�G�b��B���2Q	�h|��� ��.aP+�+�C>��V�k�+>_5�t��G!�f_������=$v��j_���-Kr,�R�XS��=,�jo�� �A��+Nt����m�%�K����Z���#�e�����W��}}��u�<{������"Ɩ�����v4� �9	�CCT���:!�߼����x��|6��"z��M����r����\���o;�`Z[���U���u-w�5u�СZ������Q�zu\L����ddG���u�@��|���R���
�j�D�5��g�91{k�/�al�b��U��=�\���[�ɿ`�=dV��cX�K:lO���Z�ë�\ę��yJF-F���c�J��KgQ�r�޽���|���"@���ڦ�U.��������>˗�|󩿜�\��Ȫ�$�(NN֔TK�I�������gF��94�S�,���*tp��aH� Óa��f%S����D���� � �z����T�>R�yc�H%P��2�x��ԥ<�GKKW�L�o΅UO����=|8zmٯ}���~���>����"5�>iT$?�=;�Ɨhk`�s3M#��荋�\_�߄g���w!���8�yQW�1@x
f�K%кs�H�M�,�L��0B�@���ƾz4���]V"[-������ZN��?��W��ϱ7��/v��Y�5]uB0�G�%uk��}����J#~�g�zb�P-�h�gVuf�Wu�˝����W��]-K�z���קD��Qi�U�*^��2MQwq�{�Y8��7	 Ua��)�Y���q�:ec��4y�xC����2�.�Wsg�o��p�w��<}ޢ����}_��~�]M/���ߗ�9 �;}����V���0B�Xڶ���Ȫ��%�Fuq�.#�ި:$�h�ͭ%��rm�v@���2h�BO.�Ǹ[cZ�J���c�+J��,���R4��z�x���Z�U���ܘ��Zgs�s��y���@,�����^�`�kT�7��*X#]�BK��5?��!��y�^�<��;��66�=�"9c����6�S�/�,xڣWˁ_Q@Y[XA��E�H�q�6��O�/�K���%&�k'
�� T�<}���}ꎺ��ܳԄ쩤�ī>��ծ���Sbb$/D�S\,W��s +-��C���tx�{q���0����B]]}Fp�ݥ�\�����A�����6%ԏ���5?�fs���ޣ��r��N�S�����slJN��+)+�c���S��7E�1ˡ�ë����pͳ�r糞�W����Z92{)��*��|�3k�4����NnI��*-Ӈ6A|�2�x���C�w�9t4 x��^�ZK�L�ۊ�n���BOu��x���cƝ>���K�j�&[$��9�g�$6@6r��_��R,R�/�)ȟu����I�-���r�!b�\����v9$4��u8��YK��x:�w����?�rc�������跡㝳r��=�d��LӞO.=�Tz������f�C�E7�����bDa�,��I2!E�yy�Zֳ�$���]����ZZ6�*D�Ti�)DpZn�M�Ն4���>[��g�35%%z�bE���_�D��X �/�.?����Oul�wG����V�b˴�Qg-^R2 a{���0�7x>����P�%8�]�.�}�TI�H�F��HFfze7H��JG����QL���7*��)x�6w���S)��h�Cn��4��u��/:w��ۖ~����,qz?|6�	"�/���:�?�"�9X�uָjo�j mjn����H=<T/�{�"89|��X���\�`N?&'�66o�^�����{rv���MC�etq�:4���8j*j������kJfU�t��d�+vv$����Q0�>7���)j�T���z��r8�'�=NX~@�ⳋ��C&�:ʥD�:՘Ca��e�ߞ����c
}33�@+{���S��찺��tߔ�u��O1]��I��0{/��Ƽ���ΰ���e�_c����'R�8�P��j���洬�&	�Q�`"H�ݯl`��~�A�t�����|,�N�9��r����
������_c.Rlu�/��JӪQQ�}K���{�'���$�����
_P�h��a�ro��}�>���N�CF|�B�� C��{���_�����{�DgM�J��jo�Y�i)|�R�������gi�"� �S�� ����~�פS.R.�8�nϗ�;}�pR�ډ]� �6��2��ӷ�}�"ovy[��e˃�lT0�I�UvAǎ6{3nx���meQ@���z|u�
$��C\���59#�\��V���v4��o���t~�XX*O�fu?x&֦�T �u����q��{U����5�	GZ1
v��Z������{?�[O�Z�O�Ԋ��WY�xO?�?K|��+�����쩼%��Ҥ:���L��Pvvvܛ�_�$����|�stp�����X;�4���&��SbB�bAsݕc�:H��%J��O�V /��S£�|Άhh��ܩ��Q�`��}A�&1�;�S�� ��n�{q�)֫����W���Gn��Ԯ�,�*
���<:!���&5���Ȣ"w�kL*�n?��l�'kN��b���	P+r��}���+G���T8iX|u���C����0^�W�mQ�ńK����Wj�K��_�S0(8{��;A������z�e?S�!���	�H�mmꗗH���xa��k�
$����a�O�S�n�G�ЖC�42�����
����vw;�Fo� SI{��Y*hȈ���4L$��s��6�����^?�ɯG�CC�nn�d���8F��� df�»��6��TӢ	h��3����WW|�V�M�2�h�
�0G�g�}v��7@�H�f8�ƒXu����5&�����~��0��pM������:�P�o8j�$_R�Z�ď�ٽ[߷C�>4����uCq�Ȣ�f��4?������P�ӷ&��4��� FKWs��~M� ��Q�$��ǔ�=�����w�3�Rq����(V}��������e�ݖ�DW7�����+���%��^�Q^p�u����� -b���`(҈�K0� S�q�b.��V<4^�m�5s����ݒ/B���R�܀7�}W|����f|��r'�8%��[�Q�xj��_���䚟����U7u+�����1V0���%zJ[z���Ŭ�������%���72V�R�1/�恊��h��*�X���{����7���ei-!�4x@`�0&��qSpg<�X�m���l_^^��:��)�m��Z�f�2� ��!�פJuA-��įr14���q� )A��'"�駏�X#j�f�[Yyx�\���������<�^{~�ͣ��^W�Y�Dy�O??;�6����H���WV���]��i.HO�������C�nğ�[ѿ��ܪn��#,ybb���x��� D��ښ�A�=]{F�D��A澎	��}2��~�S�4�d:<!��G߄×έwoO���QwZqTU)c?�L��J�kF�/����Vl���u��[�isb^�W[ٙ��tQ���xd����wԻ�c�~�-�SQ�W�4�^�yP�~|i�,�d����Ç��$�z�a��}?W�s��@�����������COKC�.8�(�����r;I2��G5����+i�_���СB��M�3��1�jC�-��T|�����<c��ub���hۆ��Yw���U8;\W���}BPv����>����O/cX�gi]�e%�r�
��TІ���_19��şs��EE����9:�����ܭӕ�Jc�0�ㄑsӐ�'Y����
"`^?���Z3�P��q�uڬ||���d���}�������B��~|�d�R�Y����K����)4ӹ0[�u��cʝ��rB�~�ܿM�&����ӈ>}{]��jGH�X��~<g���$N����p̱L�"^h\(r��.�>>�V��}����޿��i��  �Q"�������~!h'�E颔���? L'&|18�����K.ͽ*�H���m�3Ĕ��p+<?����Z|����͢J��8�4(^&��XI�'���n	�ɉ֫��e�v�HI��yJ]�j�9ƞ�^ljZLӀU��ivy�W��|���nbbr�5'��֯�L��a"��Vj����
|k �ۏaC�J�ll�����J��K��;�d*���Sr�
�|df]:�d:�t[Ƅ(^M��S�Q~Ƌ�%��x�3�K�_�d��Ƿ�?9eeK%���k�[ZOR$���ʮ`�z����ܣ�q�}��F mўA�*rZC��0$ �}S�t��=.��ĠN��5�O
X��W��ńI�=���7��i�ԃ���d<���3い ���w(ܸw�{�k������'Ζ��J%O�_?��e���P���N��'�Ǧ ���;���s��)�5Ga���*%��_��&�n�o]����@����Ss%~O�Þ`����0�5�`����}������*y�Z@Aǝ�z$\��h�hƞ�����H�\cˆ�ʵY�����=�f.�10�2==�h������h#�;������s�� W2ȉ ��gŌ�U��FʱӄP��3�����?N��{b8����h����"��:\���'���K���ޣ�ɡf� ��DS�
�T�L�8�˾������ʉ*��Z�ZUZzzay�8όh��aUX8{�C@h�\�/�KX��d�y��֡,�//��V
U`����k�ȽR�Oy,^W|\MD]gU4?Z ��ш���0?�B������!
�|�O�?�3����s����j[, ��,w�uTK��~T:�.,D:D��>��{3��x[WWW���]�Hp����+yw;M�MX���M�6�!v��������5�Gɴ�Z$0�Yv�j[��/V$2�G������ou+�Lk���
c:�`���wØŦ0���}�߹��R'�s9��y�dnJ,��a��fya�@����O�l`�H��w�:4���o���jL��d;�}tp�>�lf�L���MW;B�!&�=�٧��$&|�@�{�*ll<�Я�4���7Wwq��.p1u�����4vh�h��#x����R0�����?��i�:;_r�>���;>~atp��*Ū�B���/+�,����,��\�Ƅ>.�T�:7���y��E�g��J:������^*j�����V�d�ĳ"��8�4��ğb�w7�������1|�ňpwI*qx0��H4��mӅHfJݴ�h&�[�_��bۆR���7T:!ae�MM��GG��~���SY?��B"��]NE�	Q� kz�g{yn�x�)��uV�:�YYE
�����'_�$�'����o������J�0KQC��S��'�ŭ�'~WcS���K��q��r�Bu���x�:?02��7l[G��'P�`�=��&��ER`0�ջ�H#22���MS�;8;O��z6/�&cK�%r�˙׿����i���̅,���!R�4��� }K;���`�h����
�\� *mr�� �?�������J��!��r1 o�ӷܴ���_G�
8�o�u-|���KsB�D�	�ҹu��_��ς9Ec�d������b��jL�;O.��N?I���y����?=����n �]��r��$�g��g��z��Bv5jz�m��G�$��]�4��+�͋�z	�i�?r���7*������N/� ��T�ٹ��������z=����ٻW�|Y���#�	��O�5�x�c��3H�!�;B�v]�Qa����~�r�tx�K���}�:߸�E�np��3���iR�q�� J0Z�+o{�|.��35�O�SO�������22qn�Q-v@�:2I��i�����s��s����~�����Ch�=%�Wl��Ӿ������}���2=�?�u(�>1��k0�%L�O����;  ��z��F�P���j�����C�8�XHq{�>���3��qtU��Y8��+��+�A'��	��켼.m|WK�,yKJK��>Y�B�ዟ{�\� ��$�Ǎ-������7N	L��[�6K�`�;�Q��f2�6`	ع���v����A����t��a�/Hٱ��D=$ҧ�:�5���wP�8���̫�;�����|llF-Q���ǝ��C_��������6�.$OF����OQ,�u\����'�j�ܱKKW�mm�r��smv��2?H�w�t]�ʛ/�F�6�DC����?�z�iIu���"��Y(����/Q[��5��n���?ݔ/�H,qsbMg���u��Qৼ��-�(�ߥ���%7Imxq�{u]W��"T�������6�4uݧR!��Ζ�-saD:���/_��N����y�Ŀ��=4�S��|{��[X�Rb�/���C�����A�|'S��#���Pg�W�-mZ�U��AKO$�5s2�V7�-d�Ȁ��2��j�����32<�I������E^���!��HN<�;ې���)ڤ�d�e*3)ָz����1�dQ���00���:��Pewh�B�Y@�r1QP�2�e746&:!KKUt�3�+a(Nt�ǘ�V��a�,
D4�(���r01��5@�]Q���G�`zh�������%vY|0�{�-��r�EE��p�%���0��B?{Aף;O����W3ݪ�j�'tr?��z�5���F<�"t�ϫq"X7�4�
��o���K�.�z{I$�@��k���i�qT�k�d�������.�,�̼2��#]�?��3Y�ך,��I�}�[�3�����ۆ��βm�R2���MH;lu��Ӗ
y,_���8��U@��̀��@�Zu�������H��/�n}n�3Z�{��-G��Ӳ�xJ���Nx�Ë�����R��Pq4�~.'YnQ���넣�Qʽ}-ҟ�i�v�W�{H�#�����S�9e�h�VE�7����!]4��WjUW�]���mc���Ã.w]g�"��|дF�ږ���$"�,M8��S5�/|����s�������,����������_��B��@N���]����RJ�U�m(^�.`���~��߷�/_88 ����=�G�6�:
}�Ԧ_��-��e��I��&$'���5�_��BZ/��H�ۦKG� ��Wp����������� =$ٷ�N'��%���.0]�I�_�NOp�0�S��`X~�2�K/Thhͤ�B)��:����S��3�}1��t��vK���(�R�e�#��_[@m�~Ӯh��\����nE��+��/��Tܻ�?g+F��������N�t:����g��\(��/_h)b\�O�:>�ڡ����V`_�C�3��k?��o��ND���q�;<�ֱ�F��ڞ+�irF��z��ˬ��E�cL~)�y��	\���d@Viy`��p��=<E�b���j�}-<��e�o�/X� ���Z�E�fK�y7�p�j2��@H��
��>�rQ��>R�#��� �J�����`]�d]�U����m�*�+22n0��:�Ak�E��,�t~c����;kp0`�)�ŗ�" �hk�Jd8��2�zZ:e䦡V���Ȱ���0��+߲�<��S��w��P	��� Hem���/?������cY�Ŋ��o
Z����$t�,�,��YF\�m�I�A#�	�F�N��@?��*~�9ְ�Q�ӊ����K�:oi��]e�9��إ�zYFzK?~ժ��P��T����OO��+]ⷋ��F׵! n�rI�����M��M� �B�xjE��?������yp�uj7�blo�~��A�K2��	�̶�fW���cCS����L5�:����D��P�(E��c�:�y Ю�+ a�%>�M7�����>p��oi�ll쮭�#��$�		>���>��uK�Q�k�[�����/Q��7;e��l�V��D(WU�-
3��n��p�ĕ8�/ٿ��{���/6u�yU(�a�G��կ{X���?+��2�=�yT�;%�s�g�������Q�l�h���y��4�2&��u G���O{y����]y|�ͣ[�z`lx�8bi��SvV��ux8uY��#}曚������ͳ(;����ƿc����}yy�d�l�dS*+���n�����@�9��}�:Q�bu4���:���YC����`�(&�cWC��~u�A�����9��_<v��g�*קIV[�n%�򮑢_H�f��ߍ�u�R'2`z�k�M�}�LBU�
p�R���|� i^�(}��|�`θ�8m2�+2@nTF��2V�9%>��f�[u�a���Jm��?~0�'��@�鍩�E�{�_����{�H���-�x�d�ɩ�^��k�r�� �����q2�n�Q���NP�3Q���=���\������u-��
�n�g���O@PS�q\TA"lA����|(]��ӭh2k��Yt�	#G�󁙝�M�7�1y��Փ�w�Ybs��H@X]�8�7��Լ�[,��{6��U<ֻ�ݿ�Iq"�:}�$b��0H�k�;���G������};6�F��n^/���Y���ZY�r�S�wii�&/���ŅYT�)�0�rɓ.ZJ���F� 
(��.�߆�g+����f?�j����jɓ����6�͗�A�[t�
�u4ԿM6��Q�?:z�Ё�"p�0�:�Ѝ?��� O�"2�("Wb�~qd��˖���+D�ȧ;\�/N�8̭��1<�͍�]�-�x7c�z�<���%�L��
�:��$k$_���.Lx�$��| -��u�s�
KH��V������m��WdW����y��\Q��M&a���8J�M�l�E�;P���j['��;���O� R|}Gw�j���1���<ׂ�X�H�+�ǬhU`B�hT7��c7��χ���PH����:.����W���Ī�����869ۉTM��j�[Ȳu��<�V9��5��`�S�.[�n�-�������(@�F:���&=��¶K��tqpɢ3
��)��c����Vu�'�889e���r�>��
��� ���2"A`aQ�8Q�eD� f�k�c`|������e}�r����%�I�0:��A��&0�|�2J���zrk�^<{c���@�P�����
��I�i���[�Ӝ0E�]�x��7�*ol���H���:E4e��0�IG���+A9 ���o���b�����`ۀ;piN��P:/׀�
m���O�?�p.��R#���B��ľ��*�xW)�T E�4Ҫ.�	�]�Ks3%�B�x�M�װ�S��!5a�P�J���Q�p'T2 忬����;M>�'I�_����FSS���j��Ys�/v9 *��S<�?��	K�k�����;�Z��|�q���J:H\�#:��U��d@b� F��ʮ��T�U܂5*?~	͇�sB��;�P�tNq�]�N��n����Pͳ_���D"��`Fj�d� �ƅ�^NA��T <ew<[-^�T���ڹTB^��P�.b
? ?��q_���˃(1�j��S��r�:P�AA����`99��pn�T�[����_>��i7�_��7�ɮ�����[�����x?�`q���'����g͵�p��A|����T� Y�,]^���_����v��?n#�9hP�7y~�����i�Akc���|>
>�1��N��Z�Գ?�0�~:�\�?~���:�rr'�l���!`�s��voTq4��.~�;�npv�e���~���W`ң�C7�\&�2��l�k�_m����|;�R�� ��e���9E�S�P@����xx���Pß?#,�_��\�rܑ. ��A���^.�e8ޟ�yu�v�	���g�Q�lEm�4��o��BL�JN"����(��T7qW;��L��*.֔�/���+m)�(���ON�3����y�-�,�l�~D��* �UW��ҭx�2��ޛ�=�q7(~mT���ƏaC�Նjh����#����=�s���י.`��y�#Α�$�������}�!�v)B<��>Z 166��C&�3�Ō�ny��s���T�`xQ!�%��sO��Gǵ՞ѳ�A��[�]�@���9ܟ�����D�+q�a*�A�yM���%�l�/o,P;�rfJ���
�����B�Թ�u��a�� #X�]���6�-�g��QGy�|���c��J�Ұ�!��Yں�7gm��S�C{{~㨇#*QQ�������c������NDO�'����g�׬��C',�?�n@������^[��$�[��]�����"wi�rN����"j=��~�����nF��^�#w��e�S�Z�9]����}��Ҧܺx)�_6B���=Ju� ࢋ��q�]�B�r)w*�Y\�������5q��-.m���-w�cS�%����Z�x,į��^���LG����(
�s� �!�!d��j�h��&"#WYyӆ���B�v5��36w+�Ɇ��l�˔��K�|Q��6J@�(���/G#�;ǝ��)�e@2:�A����	rb0h�u|��=�WD�Fi����	��}hΤz����:�/q#��bJ�:df��U�t��	��Ŗi�٧LA]~!�2�W�f��}#��w*a���.��>E���L��(`f���.�	@�����V�Ւ��a����s@n����#�`��)-t��v�+yfff�9,5�F#�u�������߹߿.��vgee%�'�DC���´,�I2�8<ԓ�����vφ�5 .�G�Ã�r�s9Kܿv(�B�k��_�
�\>�6hAL���Vi�uǱfhQ�}V�i���P����Z|<��C�� u�H�F���MK��zz�b����]�ȒH�G����`��
],`w�p�r�H�x�ٷH
�{@���ׇ�4��}�|�<��d���\�P*_\��[渀]�w�ýϵ��{(,34u{����r�Ç�(u�ȥ�+X.hOf�cF�n
s��8#c�{������g�SR<��&���X<�`��nf���QۆK�Eѷ�uZA�҅A*�,Aio_	�RA*B�/����1�F���#e�s�%�+��m�
V	�Ԕ�uM����Y"A��x��0�31��5&�K�Ԫ�T��]_T�7�%(`_���5������$��JRZ:���M�S���������ͯLOߚ$U'�� 
�9	(����l���d�;	��~���vV�uJ���`B<;{&fu5����:s��\�O����C���l���E�/?^�+�Ʃ$v�VCok���Hrt�V�6�w \�q,t�Pv'-Y�_�}6�?��"��Kwɨ��8��g�	���аn����V}@�~�S�H� qy��p�kg��˃��`[�J��wyu�M��7�|�\^�r�u��P0��R��H��+�ϝ̥
wc#�k!{s���d��!���_�ږ>� ꥒ�jS�񃆴z�S��4�*���}�h�d�j�3g�J�$�����5?���z��K���.S�I�74A��j���_:��t�*U��g����n�����s0�G�l�����I��LD;��Y�x�M�����_���'�&�/Dr�.L�BL���i���ݒ�Ḧ8���IEI�Y�����[�7+$?��]���
'������m]s�|h�Ii�
@�, xcbx�ŀ}𠠸X�3M�����r������ /S�s��Z:�i(��ԡ�%�z��vz�h�@�n��s��	�rR�8A��@��ܢ�K��tt��#$�d�k*��˯��zBo�� K��'��������ᓱ�͏�>�Ք�?�pzfU�p�j��gF+�{N��5�s���+M�>�"�!|*��-�}���t���Q~�! �}��Ŷ��s��-�������x�����17�K\���ǌ���{c�9���1Tض����
 ����\�ڶ�v ���G��T�a�yaϪ��uɉ֤9ޅ�E7�.h�ŋ��Y�k�^��d�iEmUG-_�a�ܿ 8xi�6	��' r�xH7R@''eB�b� ��!��n�],��_�v	W�ԡE7�����=-�y�'�?DOׯ�x"�B2��V�,T�X�,��ӻƼL/�a�SҐK�y��ʷ�Mj �����	��d�rs�krz�)}��ٙ�Wg5��=^�W�U��
:��)����<M;�l���7���������Ҳ;��A�P��_Kl�?HU���s���`
"*��h�ZD�;�����B���o�y6LN�W0�>��4YZ1�EC�V������μ�T�.�[?���� ���ڠR5 �㮥���E�����^���>�r؍ ��>��ù��*�����v��q��:����RRj�s�1�|p��x����n���saooR;8@��.%`w�W�'�Z�,wҲ9��c���e:D.��m|}g}���Qg#�+!�n"?�q������U#ߍ��0���Sq5����?թ���v�yo�iUU��F�����Ֆ�,�rn��f{3�z\��,�<
�o�b畩'ں��� UlӒ���@~��Q�eo	A]TBr�A'*6UNf>���"m��HT��9xz���ei��~6�sH�Q��..䮮,`�Qm��]G�ބ��g)�e��U��x$Ze��<��"��ٖտ��:^sњ�Jg�_��8��:z�����>��{�z�����Z�-�c�4���+��y����	���,�LH�����ɿ��e���/?�I[��@�HgIҐq�*b%ž� ����nD�T`/���h��"W5�r�% %�NI�8�/��|l������H�x *�2[Iֆ���{3�~^�>����ȸ�#�SG�s�ŷ ,����ڒ�V�_����Z�X�p�7`'gB��TC�����l�������Vuvqc빀�[d3?�w뛚F�� Q6@������@�oj�st�$U�ht�����a�����7�@ܼ�_�8盤�Wיbm:���]i�R���R'��&"�0�gb���E�\BC~Q����H��@����g�����4�����;�����h^z�`tٝ.��+UU��c%Vu���=�>�V6�$� yn�t¶dw����/f��=%Q �����۹�o�zl՘���K(��{!�
���d����c���B���ݵ�;�nA=m,��T{%|3���/��P�j�~�Lv��݌G�}��r�1�x��P\�.��B�0T�L�'XF<�����N��p�j�p�=jѴN���'A�s��iu���n�^�I��r�[�����8�b��Z(0H��ބ��.x>��9j��Gk���E1�Z��بH��#�u��m�����A����.�bUd#1K]��b:���N�ͩ4�T?��=������FH�+ ��ۛ��{�|�Db��g�H!%<oG߭p����ݐ�������v9)M۬����}�^��eil��wVV��9���v�!hr*��,��'�3�8�0Q~��-�x��o����{�yM,�pm��K�J��N�7i-,Ĕ��=s瞧"���˖i���U ���f�S�,l�1��r�P�OF#�[(�GG��U����jsѐ��_<̿NK;շ�mc�p��1ć�bx��`��UFǂ_�'��[����0�����
�-=��_���tSZ	ݓ�ut��|yQ�����1Zn�ST?x,t�/�V?$_�``�8��Y���&�����Qq����
fhq���J��c��O��:~V��G���hR�tX��ة<ՑXċ*� 2B��!莅���! �/L��-,D�����*6��x�~!ۆ��&V�8���m0�F�D�'T�8�J#}>��f�@gX"�*-w���hhC��v��?<T7��Rb����w���J�֭� �bX���A�����b@��b*Wāg� �`)���PV�L������bz8c��۶A�����k�(OJ*5�8㩣7��/=X4�����V\����M��A��U��a� ���S�Ҫ�1��ٜ���_���s>J`x��� �Ȉ��Óv�C7�t����!X���.>/F�����%<����	��������I �� ʰp땄2��"'��ϟa�̔�m���9��B22qYYƏ���\���ڡ�K�eV�jA�<<����#���2;?~0y�=���o������ˍ�(`��a�,��$����D3��������=7���0�FH��R�g��,R�X��2��F�N\[�6�ilϥ���6p�Q(� ���\bR��g�G���8����N�J�_��{�>sf>�x��>�IT[9tt�>Y��Lm��S~�2W�>E˴�x<�$�Ѐ�H�_>�@���a�Cm��M���|6bnP1��_�F�qc��i�4������3���{�P�}	ٷ�$�dߍ5��dI�}��}��3B!��&��i��������������?Ǚ�o	s?��~^�{�{��F9�a�H���u2�n�zuȝ�����U��!r����{���O��/E�mks�7R18��+9fO��wփ�3G�}8�'v�Ν���V��r�ߤ��0-�2��*l�C��DO�������v������y��,��Q !{@�~.��g�yb:#l��~N�����м<��*sL���Je@g�7(#B�d�z�2���m)A����R��$.�P"45?�<i_IA�R� �
��~$"�\艡Ӟ�g���g�8�6b�F+��svv>n`�R(�����x~��fF~`�����6���J��M��55*d=��/�F�D^�����s���J�X���߶>�x������.�P��6.��2���Vю�Aq�#�F��t�����$~�e���,z^a���� �;4���`�̀��E��y3Q���+> ���4��NN&r�������P��.CZvq�ؠ���m��t�f�	W��FQtϸo��.ҭ6��ܙ�(l�.��0Ct	����4_G~�OYOD�)��AL�?(�&���C;}������㬷��ʚ}��{Rg���*��|����%XN莬��s����!~� ��Z��';l��7�5�9���5l��Jx��C�5F�):��J����?�\�����nDP�Y�3o7P$�e&63�HquG��
=���*U�(�.cx����k΢�a��_�$+G/��zR�d鬙�[�5``�M�\�ɕJ�W�����2Sd]�6�r���8b	�ե�8	8I�zJ&�zQX��Ǫ��t.@�Ӯ�\�y�W)V�4��������_V%�kl�R+z�w_Z[;�YM�[)j	N����O�l��q��������u��(t8\��ICE�址�?G��x	� ��l�C���Tc@̭e��}К�Tf$���q2'	ȣ�Ww���,"��2o�^��U3@AxiՇI���bH,�p�ͦ_�Y���N�S��G�����k/*[�P�va�a٨?~Yt�r���QHP��+^�	'�a񣄸e.q� ?����8Ջ|�*1��P����S�κ=�:w� ���h׮1�9?���CF1������0��+Ɛn�*+���M�(0���<���/��X�Kр�U���<��f֥?m��-��)&��� �hI�*or0��2C^4����M���q҅*W�|�!��ƫc��J�'*z)"L��$�dAZ��r�z�x�W�h�kKB{�-����,B8���ip���G� �dέ�v�@�cn^�q����ߍM��T�Ѥ��|��F�H[*�L��ϗ�Ӗ��wrm̅��nI1j��>��{�Ui����iu�<e	<
(����qޛ`�t�3�0"`V�֨�[*ՆH���ۼ����v���?oA���X��K���hdT��s:R�Y�m5��^���Q;�HP�&�e����&����(O�,:���I�����|l����Aލ^	�pF��+�-��|�7S\�hre��'����&>��=�b�a�o|���fl�)��#8�̭ˇ{��KK�7���x,��������c 9������#w�)����\/��0�M��o왛����;����L���S}ڝ bQk�8
�*�V��Sy���&�ه:�%���cs��N�"8�����@�WZ�aϔ=��q������rne��r_���mf��,���JW��٨d�
�����+���r��_�=�]W���p�_��H���E�m�O���͸w����i��͍���5;�Qndj�(�ļ�g���9?�u���d�y��W�B�������[&������H�P)KS�u|,(�E��n��ŝ��Tq#�(���T�Y�g��˖�J�~�Pv�+v���&�28Iڀ�����������1>Q2���I��lF�vg�e�g��/��C���& (]?A�bۯY��(����9<ޠ�V�B�}
�PA�H^c��M?�/�.�}z}ʨa����U�?G!�O��r|[�������J�����x��B0L�>ց��O7��~}Ɗ�=M������*����k�V��I¬eB��L
O�d�g��j����f�&fW�L�0��V��|Iq���]�C2�3<��щ�F���I�?z�_f��=U�����F��Gls?�{ʍ��|�:1�[_��|:��?�&K&���f��$�sa����ki���AU��l�}@̬ll��	!k>�..=���"o{z��x���eX}9�n4����ا��NK���b<^<?�y�!\�Il�|��5Qze�[Nɰ������F�V~��GG+���xI��ˋw��:�_i�7\U��M�d���2����3R��6��:����n��b�Q\���2����<3ޘ=�R=��,n�UO��9�~����% ���

]�G�G4�7$���1+|�ӝO����ϡ�n��?X^]MG�r�s�Tg��^eX��鍻���Dn2�_Xș���� EEDF0O9��vv.;4�>IF�B��wxb�L�� ��  �'����F)hg��,�.mX�z!��I�4N���_*ֻV���L�ĸ4��%�Y�����~�O��{-%>�d7qB �n�n����̔G����yw�rM��Q�H��*��ȝ�*�'Ԓ��{�N������';���߼����ki-|K7SX�9,-���5�qz�f���j��L����ןk|����,��#^��6UcA�U�{p��������8_�bI��x�q����Ĭ'{!E�:BO���h������X�;ifh�T�^P���r-@�`R�0@�����P� 
E��A�:*`W�f݈�����������q14L�~��K�v�mr�����@5k�A���k�L���U�?{��O�\��ӧO�i�:�7�^W�E``*��о��q0��7���5��G^�R4��]~���<M��=�v*���|�.�n$�p[����ёn©5�8�֭[��ƝD����<��<��YYY�r���c�P�uq9Ǟ�_�d R1N�H������CA]�цx����8��gN��/�S0!�OL��N�
֑��#O�����֠Ő�S����ư�z���Iɨk���k><y��/�$u+2g=Z��M\���߶�c���w��)�w%S�u*r�iK�/��]S�u��4���pټ�Qh<[k�l}�����8®;i��2M��~�4rdD��,	\�hN�ʰ
:����C pN`�hI��vt�C�	^W&��hGt]L�Ҽ�~��gda��0��x0����ٸ'Z�S}���^f����z����D�Ѥ���K)>�.(����㮆����
���T����م��c�i@��	d��[�7��~5l������)��-
�01k��'<�Ȉ�i�W�K�Ҋ���O
-Ԕ������XԒ'�n���O G���Rl�g $4,�O�@�_����_�*�#` Ύ�4�#W5���[[%�R���U��
*T�fv�%�_��/w����{��� >Ç1v#��Im7h�[�J���%ǯ����PV��]ҫ��[[[s��cO罂.���5�?1311�m� ��p�� @eKKO�����Z2�(A;�S�ƈ�Z�w��m[�v���NQuړ+�/u`�/�B*�k���8��㓗:��4�'�����-��!/ߤ��(M
����z�㔥�FX�o7�T3��@�_Ph�'s�%�!�om��Dc�@�C��ǫCv���a�{��`p��f-�CI))���M��Xz���p�v�rr�"�K�P7x�����p}/��5�����A|S�",��W�Kn�r5����)�r#��������`f7-q!`'i�LAwx a:k��o��C�i��L��l����z��S�pT_�����0>9��,n�߃V��2��S��3�=�f6by�M�o�ђ��MW��U�B���F����w&7L-,���
й��4{�w����t��YnKQ)q����ܦ��@}�ucB�-4�i�E�z�����CQ�^O�A)��	�ؼ��$5ogIiZ�~���J�*$$�t��U�cwwR����Ζ����ww��p�}����c���12q.�uΣUXT�Ġ]@F$����as�T�F�W�H�)��:	~2�B� �'��i\".�+���ٓ+�n{w#8�o���MO&$�*2�L�W���n>�!�[Vl${B[�<�U�|Z�5BQmH�DYg4���Y5���(�&ի�0}eѼ�m���C�rq�̀NP�%eȁ����In�\𰴱����b�r%zw\)w𽥯/##����իm��m--Q z7��P�FFʠ�������/-1 ����1� �A	��V��3�P}����� q_{�xf|\L�* �@6���ai�y�s@�}�3�W�3�$G�+�=�����9�	v�'>-2��eF�D^�.)?{b�K�R���~Y�U����JMtag'i�zkϲ� � 
I�"��� 	!(��d��N���̔���OL\�7�F/m�m�.}�O�I�FI��3���񀬜����PY��r��-���
iS3t���������������SV)��A�i߿ߖ���I"6�d�D-[9����Q��[�u7i,�������mb AP
ޑ�� A��5��/(p�����U��qe����/{����PFb1���s?á�3��逪?B3�ܚ�q���E�@΀a��� �dSK,ȭ�ͨA�YB�I���N�JI
0�~�.�q���4D����l�.��7��GC�5�构�zɏ.o=�>@����R�	~��s7���_�9�i ��Q�6�Wid�\����нw|R��:ghk�$0��@&=T^Mhj�$1s�f` � %Hv|��WfN�o�:��qc�8P��O*�\*��%<1�zh�-��K/((���摲������O
JJװ��l{���X�����P��M_6���o~V�H����B�9t��N tѹ��R��,^�z��Eo P E���׫�dA �ܞ�j�0��C�S�����q�ěb���2{�A ��L
���>uj��;L�l�n���?ܪ�����N@w%�h{�%l.֔�"���Qc:������TT\��X�U�	���m���<�e�fw%�I������JL�c (��M�@�ʿsA�=����婱�@����(���V�M---�zx����� %�Qkj�6��)����۶��U?��d��ٌ4�yAS7�ɑ◕7g�j��Ah��]����X_w������EՈu*l�%��efC<}�"�����:��w���Ia�DYY�/PlX�����/����*�檝澜\2���|���e._���Ù����@�\�Y*�TV�f��{-GLx��c�/f�_�ǵ�߉A�[[�X[D-�:������	ڧk�[�N.5[����屛�+w��x���[^��Z_ y`@��;6�"�9���P��X�i�����޹�^�Δ[:��ikO?�C�2������3a��U?�*�,�r���܆�Ā�M��ųC,J�T���л����}�����_�R��J�)�G]�N#�'q~��G\�<���ee�j�Q���@فcR*�y?1qh����4;��q���91��S!���Ԙ���j屷dd�US�y�/�d�;4&4�[��� ���=pۮ��d�x,p�X{����OBg'S����+#�������	,VA4��ZV�|��bMq5H6��D)VSKC|��,ѭ�4��u��'{��I��.�%L�֚<ƨCo=��E8�����gD�Jc+'�)�^�6���T�繆B�\(׮��ރW��ȃ�TF�LS��� +�T(�m��q���˓1 ���V1e5Y�x�)���Y�����,	�q�:͑��+)!��%}��<?ur�����Ⱦkn�A,A�7���keee4��������P�4\aec�9�ǣ_uYȎW@���P�ںW�}�����v_�v�$���1o[ZF0�z�Ӭ�GG� -�т�u�ϣ޾>I�X�Aw<���&gc��� ��(����?�(Y�Ir�l�ԟ H	���NQ��bQ�wɑ��٧�|�ɒz�p,7@<Cΐ|�w)�S5�TT�:����/�˃~�z��I9���À����A>WU]��6'&�+�3M>]=������ ,[Z�c���׳��>�
�W�.|�����	��|�DG� �
���nI�;H���Y�
ޱ� �k4����oq�D5������/��lF��7n����y��;�oT{�T�;:"��weUS��ۜ�g����յؤZ�Y�l?�����5D�Ԕ3�z�z44I�Z^�Q.����hdUu3O{���7t�	�Uڳӱ���q�����33����9����Ch�i��[eƜD9Q����V�E߼٢١j��J �m�v!�>�����?}X02S+Y�1���w�)(���=�1�����/.�WQQ���g�$�;h�������ttt 7z?}��A%�	i�c��\�ʾ^b$� $��n�}�10���b����Fbe�}��:�%*] 5@
_��d���oX'�'�~?G�b���֖���G�9����&&`OeN� ������L}�ߏ@�3_Dw��앍�N�´�C�`�>/���s&
'�(��+|�/��~�����>i�J	G�zhJg� @�Fi��ç}^�L�n[���:B�:��4��Όb�I11����z�£�r�vP?���������/z����˗���oyv"��e��H��-�����ݟ��8�U5���W������=E%�l�?xfׯ_oJ,	�FYY[�U30L�' ����ٹT
�Z��k�Yu��9IEwVY>}JVf/���%�ܛ�����Y�����4N66oJ�����nY`hN��'�t�z���<{"Q,�?�R���,�"�,���25͗���E�hej\%��z$���'�G9/5L��J���Z\g���$?/�|"�2�tc��Ia6&L�7B��n��}i����)iz�H!���$��o�K��_��/�p����8�:"�t'J�K-=�?�ɒ	D����{��/Ez��g��-7����9ڟ�f()��蟞fO��qE=N�<��GX;��MM��v���;u��
{�������T���]ts���ѭP��v��\�E�֭���a��l�&�{	ż���
+���&��{D�9�nf�y�k�s�en�,L�E��3�S���s�b��{Xl�,pY��Ҥs��.m��)!A�}�
p�غO\��h�;�M��Õ�� �;��+��Y��L 9��u@t˔P�����ם	�8� &$��>R��s|=|DB���R8���cMMMnVJ����
�����6��n�޽S5�ˉ>6<E��5А�Xd�����������7=�GX�ˎ�U��3�*��²�.�|���
)�;E%$�m<>՗�tuI����G�(�0�b[*�x��,��8ċQ��T�$e��fg�H�p�^�a��a+�74��PIR���2e������g��
Nj�K.	�*֠�t�N����1^�)/ϝ&�h� ���ŻȒ���+��󶈳v�ۊ�r��y��˗z?��Xs4/���Ϸ6\������-�mv����ۤ�laЀ;�\.�п�'^V�TXR2Fg�%A���������,�O�;�
=ۧ�G�w~}TЙ�W�qw,����#B�[8�M��8汱1�ZO.��K�����|����Ǟ��E�@a11���vO�&��Ǳ�����p8��A"SCm���	�H�*�~�S�)�@���ރ��f����D���+N����q���w�`��U�w�N~��f���gY�Wp��>B�B?锉��Gwg��̠�S^��<)��~�hӉ��09H�_�6��uv�N)�����<�<��k2�٨���K�A)dN�k'Y�� u�`oY�����x�_��l��1�H]������Q������|�DP֭��������e�iS�n��574$��<��jo�����e�Y1sXz�W�	S�Mm$5�T4�BЬ��RH7pV;S=6���'{p=��q��(���b�C�u�D�g'��I�Ɨ�i���?����^�K���<�0� �c�u:��& '��T�4��i�����EyʏV�I��<��
��v&y���/mA��w��}� �QH�ڻ�-�'��S�~���\J��}��	�̈�ժ�"�AG �k�K�q����4y��[=}��8��]���(�}m�����]�ٍF�����x����A���_º��$��RЌ��`h�D���� ��O�pI����$^�*��R[x1�7z5=2V��v�O�f��<�8D��������K�dsц'��4��>�u��[�w����쪪{~���J������V�r�!��v*��Q0�P��7�F-�O�%V��L�����~/H6fXի�śW�
&66hrds��ʇ���QP��67'BW�9t��̸�O���V�3��N�4�56�WU��cJ
���o��I���ww�+�	v	
",)�n�ޘ����&��� x��)��?�K����ۺ�ip^������������ʺ'm58�[�]6��k��P.�!`]b���D�z'��b^6��,o Q���A	N�$127�s�Ӣst���F��'=~Z�aX=^�n�/�����[-k�������D�\i�\!��:���&%kS�����&ʲE���R��3�p_��&7�F�������?�:͕�2zvv.�V ��UnII�V�Z�:\~��N���"9)������a�/,���	���{������ҫ�kl4��J������lp#U�$͘��mr�C�лP��A>���6���"�cx��Z�OkclH��{�\�deto��`}kկ-h�C]7���9yvu5=c���=3*`ht�{��� <���QB١1�Hp���'�<7�j�NT�{���M�a��Lh"x7P<<�3���в�X`�"�6�S����U�WQ9#�5�c��8)�aHD�v��3}@�1��
�e�J��ױ�#>��!׳��f-�g�h L��XW�_�s�β��ols����̱�v��q߷o	k;a�/0�hy®k�.G:j\\��o\��>�1$b��uo����3gPU�l��?DyvPv�}o�%S��ۮC�yW�4��Yݛ�ݘ��ȝ��X�����i([|��|�d��e��@,(I�߻�']���/EK�$���� �_0f�Lɔ󵇎8����e��-I�<�m8�"�J����L�ͮEG.z�wWwL�
!�_����ʘ�}����i����_$�HS�
	).����xK7������ʼ��yt8F�7���S&�ir�v���7  ��i0���z��B���W�R��)P��r��'t�̅�x?� ��-�w�V���8�����!V��3r�r�k�@
�'.��0��b���0���DDl��1k>��2e8f�+8Q�Z�w���n� f&��߅�M�(=���(��$"��b���IS֎_T�~Y)`!�UK����O����}�f�Ď���b�2Q��p�	��a��k�ݶ�A�u�OwyL@2���EQ�4��>@?��|�ዏWOJ1��%�ݘ����C8�fi �<���_I,O���Ɉ�?�
���3��|�+�ZΆ�����W�>)����
=^���0<�NT/��k/��9B�΍:��o�C�¨���@���!�Q�Pj]�,����D`0?���2�弲�ȝ\q���q�����@
�lT2@8w��]����ZtWJ�h<HK�⥞POE `$���^�ٴ�NL@�6����F)�֜��8���67�'Ǭ�VJ��[�Db�ЌR�|�<�����ӹ�,����7��F[#z��;���I<����`�������N
���kjn��z"�AM<(2H��9 յ�f�~㓋�e���wZtg�/�ҫ6ܜO��s��[���?��O�VA�I5��B:��򼴽ssz��d�M��8yt����G�#:��b�/��???���V��k�|��;��no��P`J�=uu��n��"dɣ���X���}�+��X�O6�+U_�}�����$$*ob�	sMq����k3B"��1���]��PW�Z�re��h�F�_ �.�C�`����f��?>����+��������)0��w�=g�.|6%a-��m0�v62	���!dʺ�8�Ā�9�zZ�/��*�ck�d2��҅�?|�J�+b�t�ɥ)L~1]�&����V^^�S��_�6KUz�����_/�	�s��l������u>��7:�9�Q�a:��⩁^>h�ԇ�^�d𗾷�"�o{[����/�m�/(���Z i$��݈�g`�a�ꪣ��J`��ǋ/8��YՕ����6�6�P�>��ݧd�Y��i����ĉ�@Uox��5�sz@���Eb(�3(��N�e:��k�5�}|������� w�D�)K��gd��Y�Xc�����NO
��K��|��ȸ-�=z����c	����-�T�f�w,VY({��6bD\��u��֏����%z�ּ4��ڵb����������<�`z`趯��w&�	 x�!���z�py@��Y�9�T4�wz�2�t�ui��\,nG��E��⫍�~G��~���j�)5�̳S�̄��ϸ����f�߂gO���1R�O�b?��'B�䪁�i^�{{A-�+M�%3dӀ�I���=x���}��xeۭ_����a��_�7��$��cd\�$�r�LCe����@\�\sH��e���ݶ���;q�܃t��5�4G�"���P�jC((`�t��^gN����n���T�A��ȟ�m��ίc��y�ɍ�#d���ji��w����=!o;:"�x�3Po[[�u��J�S�@�n���?=��w��I2v�ı�zF�;�0a'Х'����JJ3u�=��M��>��@Մn�d�P6��v�&mƶ��?�����˹[��>E�IV��_l��]�?��o�M5���hB!%����Gy�j�.�[��s�MN�8"�~��;�n��G�>�!�I-nτnu>�ݵ<�� ���|i�]��~G{�}}}�;- ���n�,]-	�۽u�(�:9�	�ek2��e�=�p�v����#`GF����O0�kB�P�ݙӫ�9�;����B,ڧ���+[�k�K_K�T�¯B�Y�0���M�c,ޛ���ZA1k����Tv��#��~��aPe�r�0�u�_ۛz;����5o���}����& �k�����Ǉm?�΍���i1�1WU�=PĖ�RP4�m ׍B/E��N���d�zU) �6�7��J	�O��z��~,$���ݗ�&��r�O��C0w�-�N�~��аKA��ݛ;���=O���s](�l&x�vk-22���S�o!tqf˻f���� �.��Q$��uu68��$��"Z�I8�H�}"�M k7�n�8 �Ȍ����	�A7y?|�4՝�d�H�ts�c���M?a)�T���� ����]0�?�N���C ��D��C#s��h�z��9�����S�q\4z)DN�<������ez�q]�l]�i �*���__$NJI���V�MaB4����ؘ?8�L�x]r����ɚJ��1��Z�gI]c_�8���v�{Fed�R�"���Ԍ�2QW�3f���8�����а�yrF�|����I����yYHy�y�A��+��;�Nn���}q�ps��&	������7J����L�~<�/r�b��U�Qss�Ǯ�T��S҈��:w鐣_�b;"Z�<1Ֆ�+I����J	}�_B�onK�l`މ��H�����ye�*%�>y��h�O�'K�'��]<���iexj>'hvY�n�h�<u�'@дw��K�0^CC��~����>�S�?�/WUU�w��-��{�N��,�� �T�����Љ�����/���d� F�2.�}�qnƞ�܁"�u6��a[ޯszS�d����:����`�x7��z�0
����^Ͳ�9�����@��v#�\HD|�@��vs{;� �	�kqqqv' �&_dd��;��Ufi����n0O��[܏�>~�ذ����d��.M�0J��o2O��d�*����_5J5�[̢�Ǫ� �+M���ݻ�U�u���J��&�>�Xizv��g;vJ�3�8nݪ�b�($D��J�yZG{�T�8�z�y�-��?��QLw�.A�쪲�%�0����4�\�9*U;��b
���"��B�њ�b�A�q��^��Z�G_74��$�jKL��R�71��M
8��B�� ��Y�M��������F=���괅��1��i�dj�뺻S�D�Km��Z�Q�\Q��đ\đ
�Z����\�}�3�`R]|���>�Y���h:v-������F<b�R�n��}���gX6
�~����;HA-|���Tm�?c�qh�R��
������W^������E@�I]Y�˛g��9���UU���_�ih�T+��uT�Z����O��,,��i�A�=d���Ƃ��o��{��j��� yz�}����D�"Wc |0��
��������������w8��������3+/�F�.Բ��zS��s���#J��%#Cf��"����Wm*��y�v���3A�.ǹ8�5���貆�)�X��ܱɰ�rۿ�|HT�Q�M����
��������!���MX�k, ^y�M�/�L�����`l�\����v�E��.{Ab�k>_��/���0����%>�Bݤ��uv������"/�
 �FԀ:y�#G��v'A���"����s?�}���Q��*Wc��u�YN�WK���R����xQQa���d2�ځl&�T&��P�<�k�{9��򧒅#�|���k���Pκ�2L}`p��0��B= (�P����Z������M����*9��-�ƵQ�
>�k����MQf�ܱ����u��d��'i����iw�`��J���b3W����iAa��.cy#�UJ��5�^��P���x�˴�H [��KXBDE�ތ�<�J�$d�ݧKmFj�N e����,�A�('�������_)�<	��!U���w����~nKe$�����Yc X�h%���7iO�U�E�%��-W|��r�.���#�`I�#y����g~�{{Cg��ꥱ)P�}�.B�c׀whh*Ѣ��z�)%��?r�0�ڲ#�'*@����)����0�
��p��E�p�ף�����ax�(��P�1�NA�aU��)̸o�����׺��h}|}[^�:w�����d��[��2�M�:#/�+Sѳ�4�d��=׸���:ć�C�5$����gO�&>R�]E���e=���[��f���8x�a����P�3
=�E��G�ȑ-S�5��hR�7��ӝAQ䫟H"�M�I��7��\�G��z�nPQ�ç�d�i&z�mc/�3>&rK�ӲE����y��X>����)ӄts���D��u�sH�߯-������v�8� �:W���W�.��j�ta�K�oe���0 �  o)'1Y�fFV5_�s�?�y����og5�u������!!=M.���9H���'���l�eݎ��<k���U�3�	3��\�����w�$B�Te��c9N��~|Zsi:!0p����9)����N��x{��2�ǫ�����_��d��! � )B���@���/������3�Q�V�m��q�!a��5QkiM8 3�\_��ˁ���"�LM#x�c��==3���.&��|���(|����]g��r�9�]��Z7�
�S���/�6a�N�Τ��LO���1r��.�\�%�z��L��fl ��wl,F��5]�>3x�M��rWUM
�%y��Sg�W�����d�O��:���	c���E@q�T�in���K��&�~��?~��k (�Om%��sˊ'�^b��u�	��{	,��?IvL�G+���pn�������a:V�����K�<��5��.�X1����Kj�s��]���󚚙�f�+^? #C;ό������?�z���L�����J���2���͒����E~v<*Q) !�	�#�h����utX=�֟p��iuˡ5@ii�G�>>	H$�EZ��Ť�Ěm4K㪓ӛM�5�m��ý=q��}�l����T�������o��v�Bv:��Na�P�:�xŴ�[u�;���3W�EP�_����pJ��~�9��X�Fw"��藍a�Ǭ���&�Ĥ�����%�?'�Tֶ�ce��I��^ON��{�av{[�����'���5�Ӯ�ڒz���	$��h=��M͍p����������2����ne��]�vr�ů�Z�v�~�,��w?����q�*'D�K`�mm�̸�si�YL[��ͽJ���̻#<BN����`	�
?Wpf��D��|P~��N�a"��-��n�V@'��5��[7!��ϳڝ������4���J{f@� �ـ.D���j�&g��n����&VU��,�F�g��ݴ����0.�r�xH"\rm��[m�d�y�a�G�����C-��q���ݑ��7���YXx�.{X�źZ|X�wq��E�#_�n������/�_G�����U�ۀ�~`�(��.��蜎���1Κ��4���x*�T�:]Ġ6������<�,k�kq���$��P�l	q��OB�e�|JnFh儓��k���4{���VJv||\��mk�3@����WV�A�?ceZZ��m�ԎCk���B���W�]O=@Y���t�1>)��uHt�R�_b,z�.�L�C|�r)�����9����gɄz*���8y�x�W;V�P/G@X8y�~��c��rJ�<?������2��n7���d;c�2)�H����@|.�W	��#��\�۾�t�4�D�:ĕ���;m��}�a�b܏�Ird�%SQȘ�1r��(8���Iw)0!�P\�9���e궡�5*��9''#ּi._u��z�y��P6�~HDY��\Dv��3s�_�Y]M�4M��
;�?�P�V���M	F�]�*��g�խ^��1׶��5A�������8Ug���I�ŷM5浳;8�b�|5I��~�?��Sp;�c��_���^j��K�F�Ts<�6|�܌Zd�v^����o��3���:�n�e� ���HЋ��"I_ 9'g"%k`�{p \|.��r�Z:�g8�Vˈ���ρ4�=�Z�Q�/$>>9�b��v�]�	N�02�	H��������,g!�1�� ��\�%�i �T�ù���^M��SS#Ħ��#��\���-9��A�2��5ZM#�cE���/����� �Kb�8�69ф��+�nL���GF٨d�? �*ȇ�XC�|ӏ01�GJ������I����b�<3	Pf�����|�--�ͺ}l����N�-��G��VU�
������F��+&��ԙr뙶����s�*
���3q��Pc,;�NcQ����㖧�5�Hd����M-��k�����Tb�kMo����i�	�i)s=Z��:�]W�ެ�e�C#����k��Ϲ9B������+"��E�Tо7�y規U�ZFOO��A^U��:Uu���(��<N���MR��`����_��¬��?!_�~�lV���n�����1�����؅�X�s����L�?���+�7E��O����?�GN��7g5�X%BSq#Z�����p�o��Hn琋$F���|B�;
i��2��qNG��:x���!v�.�ʤJJ׀.��Q<%ԛ��E�x|�|��N�H�%��Ӧ���%EH��T���Ta11 S�7�Ą�n�X>}z�ڰ�����+���>�3N�uMM��ޜ�Ԧ��(o����l����-�}6�a��';����j	P1Z[[�e��70�b�f3g��v��:9҈Ny����?I2]1@�X����L�?���������9K]�gH��Ot����Ψ!@Fn�x"���A?M�����q�f���'Ͻ��|lcC��x�/�������m����)�ay�Ӄ��6��H��/+ �֫�R�IV!rt�m�"�F�
~Se�	���.Tڽ� yI��om�/8�zn�]E��C�����(o*��;k�9;���@>��G8)��hh��w��[V�]�����Q��HUV"�k��`�U�O������iNU"yZ��Q�Dpr���CVIf>;0h5U�V�~g�i��K�K\�}�[3��]����m��i�-c��Eؓ�LQF��f��oQ;����AJ��Aj�|�߿�xN������"ŉ1)�m4(�[Ԓ3��Cx��8H�����
'q��g-�	���OAV��Ul�pE�ab�5�K�,[�48%���و���H==�N$@!S�,\�M	?�~>^?��n�Euiv��?g`@w��~/:�8�+uU��d�V�4��D>u�	�o^F�LM5�7A!!l�X�~��ۮ��Gk����s���# ��P��bY4�����Smp��g��4yU��]Oy*������(f]�{m5����ed����2-����u�z6*N�:�.��t��p^3�Q�n�^�3����.7VS[��{@vS!�45��W��}��,��)����o7 �9�z	��,,ϖ#�����[ҡ]Q��U��_��f��b\@6���*�F&���⒓���Y�#8��H|�}����������˰��/�zQg�'� �b±�ҕ񂢢P��[�ǌ@�f��w�7'ɇ��~�6x,�T�F�&���n�z��<��	 �+f=��5H}7O���y�R���Yuq���ܖ�ְ[pp�Cc���8K*�'ɩ\�/-��tY�q������7Ƈ�>h��s1�ӈ�l"�(H��R|��{�󳡶k�)�3ѕ��-���_i�bƁu	6�o����Ʈ�o�VlUlnݹݰ�������������T7�$}�KS.�;�q����S`4�˒�C-�ZZ[�zzdѺ�OM���g��3�D/y���������@:`��]�޵�����|�������M�?D���x�>|$�;��r(�������M��7���B��	�Ma��Б�����5I���ֻ�l�-E��[�t�-����Io �G+���?���KM���0����r�bx���Ðh���8�OK���JԿ:������^��D��ΑDx=��%�$� ?9��W�E^^���H��,�U�D\]��I���XZL���l���P����<x��EQ���8���v$�5���c˞��G{�D	�Bs�̌��$��t���Cg-:�'�����$�w�������1��(�@<$,��S�4:�H��O��'v�V�=sB/��p���,�p��L� N��#k>@E�h��j���sH޳�wN��D+�R��	A@P�.���Bж�5���?�a���r�hZZ[�a��mTU�荥��3��V���&q���sgr��~��7��\�K�X#33�cV�E{��]c��U�*�b͚�O._:t���@��������}��f��2{h�ÿ���Xk|��<��z�t�ʁ)O�s��EV6*n��<A����W7O�AQ�-�����gc�܌U.�@������/�"t��"�|M�Hq���	t�����;�����U���{%$I�$3\3#��M���2CٲB!d%d�nH>�n�^)ܐ������;���sΧ�_���1������Q���5�!�ӿDI�k��(�<�u�l%{dR�@�k wv��e�,�y�|�Gmln�9K��#���ё?�9��V�G�.J$�;#�����N �U��	 50�x�93oؿ�Y^S��1����O�9������ݜG�P�z�V�CxK����%؞�-����Ѿ�cI��II���'��� �8}t�r��Aj
����p �g�cZ�A�J���봵�',�%"ۏ2���4:6��4�?h�w���!���U��+��:�*|��o�d�~z�|wbU �};$9�t6n��������O�Ngo��N�����E��M�������&�r��d4Wrӯ;)���n	�R�Q(m�;��ڴ�K{�a瑱<�g~�*+,�>!�u�.|���0�b�`��B��C�m�dzd�`j�<��9�om��w3;�xbbW��]f��T����g�i�J|��)�B�L�@��1���8�'ov�l nq�4�g/85�B��Me_�R?�9.���7�i�fp�Ε}���<�mNW���-2�Q?1��n�)��������w�y�� ]m^^^R3�\��H���0���>��`�}u%���ekP�!�R�Ӗx���|��o�$l?a�� ���m"{?
�ݤ.7`���+W�"/�XqՇr
t@�qS�n���,�7z��2�5���*�3�  M���u�G�z=$��g��vg�Hv���c�a� ��O�<���T"22!����ܾ[( �0��g���֯���D.[��ȷ�W��buea ���a.bktG8��ݽ�A�
�@���1jd��6MmJ��{����hpe���dʒN�C���Ы�b�F:ѫዪ9fyvF�Ȭi�ɷ�	 ��֭���Ȝ�)�??�<������uq�u�����m?�^�����G�W$��~�=�v�UM�*�#--e��v�����~�_,Sc����,K{]�E��nD7
u]����;�I2v��%�eNO����� &x|\8�P�vv����I,rqwl���E*?9�6Y�� 0TS��Ҹ<�&S��I�Ɠ 0r�sH�gyJfv���,�e#����;&��X��eȠ7��agdp~�r,1$,�Z�W�߀!��WU�kϬ��:�I�Sn�؂�4����ME�$��Z�|dZ��rK�~wãQ ��$�yZ��������\TX2�.�X�:/���I �8ھ��G��W&�N�:/.5+���v�oo�H�\zK�^J�y��h~B�ϟ?5q�{��dh���K�o���������aQn!U�4B+���_=�+��U=����9����EHkF�*�ٞr��\��KO��1���_ݏ>�SnS �v��\�0J�R��"E*�o?H**x��������?�E5��S��!�M~�#�$;3���g�����L�6� �������ָ�g�8�ƆG'�?��0̦��k�F�7:��i̡OCBdt����U�SX�����N=9
KWu���P�e��m��P΍��%�w��׌����:�~K�LI����g������x��y&Ck�yt�}�0ir��Se�׺��Uޫ�	b,��w�1{�����nJ��k8��J�}�k�gC�5�﫾S��k����H��p�W�[�(�F�������~�� U���!��۪��J�Փ���x�v�c��s�l������Lul�g ���N֌`+ߌ,�;;w��D=ԽLɕ������j#ɦJ���_���m{%,��޺��8�	|b�j�9��^F�l0b����|�y0��H�V"�-]�N=t�t<�� �^�-]�P��T��,Sߥ�kM���F�ǯQ����=�Γ���D�mZ�R�L�z�J�RZ
��/LDq����}*�ぶh�������9���N��m���/@�T�We����"/������@N(����Ҳ���>��l��y��X=���tɓ�x� �'�))���8� �{�G��4��q���l[�A��)y��̾��A�ZW>�XH���EA�$/���R-��X툚�1�����l��l� ������s�f�0�L2��� "�K�4_G�P�;:׌ � ���T�{z/�����n��_��֮=��i5>`5_�{q���g١�Hp���ל�V�76{�����ɞ$yf^9ՌT*�<k)�ci����ǓZ�9M,���^/9���x7�@`C�fc� )ҙmiiɜ�>f�c�e9Q���؂��/	�gh"�����D5�qZ�&7O�q_Oxl-aS��k���f ����oO/��{s���$����� �<�T��mdnęH����BNv	�
�?�����}�j�N�404l�ￒ<��v߼{�	,��R��*��;���1Tw��B��W5��O����c��,�o��u)n�z�:s�F��^�{cN�ڄ�����u�@�F� �2s�K�LW��d���*�9;XI. �*�1��/�W� �m-�<n��%4���H[˦)^5�r�w�ܚ�����(�fg?�M���!N�1�/���v �>���B^����d}&߽�$������6ֲ�u��:5G��� �n�%e\�+�"P�y��vوt��/\-��*�0�6��Izzy}�wwD4�R�%:��RRR�<}A�F��L�g'�y�c��4��Ȝ-�P��q�<>h�
w^�y�_�;_��]Mu�`�����uk�YRz�4�\V�"�������S!�W�2{T��ru:{zȁƎ�Oĸ��wς P�����_���G֢�����'��gs��Ą���	������y>�Oy�>�lV9�aLxc�SG��u��mEE��~�����(t����#c�|7�{��	� �JC�#�����}ԉn�/�JA��DN�����JI4�W(����c��A�OO����ڱ�L�)�'
�ؔ�g�`���jӧ�T5��x,�PW�aLŲXǊ�m4]��uD�9� p��[�٦������Y�l�ҿ�* 4�A^A�:.51m\���T��O�)�V��YZz���z�-�Nك�}���[4X,6��LJj��S�����扷��6;w���83�I)�Ǔ Z�[Qt.rGc9F �輦�HA�J��n���B���/"d��+!JR5����ࠟEȜ�e���)�ˋ������H����#5�m��LL:eY΄�A�zIf��&��2~���������k��*S����CBv�����6�o���A�N���N$ob�Ջ�����������j�'�����s���<d��X��s7���S0�E_2L��^�}��GF����w���u��^�xWT8Hh�L�+�ã�����F�~��D�r\�o�6�t�b�D��٢'�����w+(��|�^�G��~�X$��a{|�G��*ێ�ﶴ[���p�<W�2�D8zE���� ]�a���婀�`��b�>
���*�V�Y\������\�o�r�����x��w����NMq{=g}���#%>ʧGBAAQ{#�V���s�t���ŋ_7L��i;W0��?{n��|䴜(�������2]{{/c�x�*��s���C�/Gy�A����%�Jj��3f�ra�ü3�Cn���V�sTT�Ѩ���4K#�q����l�P��e�e���1��s�F���U��9F��ϻ�xn�\��|@-$�vB5~����}x C�a����b�,,��e��m�KR�(�*���646~X\�!�m�c�䔽l�5gZjc�㫏}�r߻Շ����y��x�O�"�Q��H�'�]�ep�x`�k
9��������������U���y<�4��Ī�1��Ҧ�,�I7&�J ���}+��s�ė���Ռ��4�[�� �v�[���d��9i�̹&ɋ�|��TȻ�s�K���b���R*X���265%��?Kw��ʊ6G m����o烠kD����y7��y�#R�is�o`v�ɼ?�a�a��a�<�I|��L����8��r��)@f �j�'4�%���+�����o@?D5#ǲz�Roƕ.JI�ț̬x������<S�`��D�w���5.�9�z9ǜ.�l���r�8RIpf�B�������������N�����	�~��͸��ѿ��UUc�>_c+�ȴ���;�-
5}���EϷ�4o�WWF��>���<�H�[���uO�I��n8К��h��SBʿh��o�9�v�5h��?>M��/���?�\<�p���/�k���m����d}5C������k�^s!F�$����0+�T�'�}.]�|�E�~q�g�̟���h:�@ٰ�*���5_�(cQ�f���d!Q��8MM+����C��^��E�q��&���5fw�\n	һz{�*�Y9yx�]k}�������zڅ��ׁ�Y�����+%��9q���A:g��e���e��Z�W�a��b隠��E�W~�YK"=A�_� �s)���e���nRbG �[8��)4�]�9 �x׏��F�TR�ޓ�^��QCJ��T_$/��6²			�{x�#m�d�\Q���������U���/�C���]H;�ݩ�##S��*��-�B��>8_߆�=��66���ؼ�j�yyr�K=��ov���9^��9Q��=�_��i����ν)�Du*U��"� CT�U�2E��J(���E��2�ْ9���=�-s�N��b{j��i��H�B�
nn����+f�sK����4װ����#�����-�QQ�߽���e[�ջ���S�k.�����T�enl�tv��Q�� ��:��-��8`~���͜�������y7�������%���A��6��*�=+e�W�0�6�Ry���e��>�>=�8����0��kb���[�QiЖ�Z��6*EF���}����C���PG�;nnoj�&=
V=S.��1�z�Ї��{�ccn��Ky�"��eqӝ��?c���� ��=�8�B�[���i�zԽ�݌vـ�G8\����g/��H��殦�Ȣ�x�.G)��˽��֚���yԁVA�r��el�6K@M]�DĮ��[�8�u���9�Z�����]M�]�2fBY	���Kӕ��nm�9�ėX}�}�:��af3���U���8�2���j�VH;D�zg�1$�I���A���ʥ�OF/��ܢQҡ�@#����i��(�4�M�9^�4H/��Q7[�X]$�!U�n��gLĢ$n��ܹ&ԝ� ��t�jgz�[��ϟ�yIxU�\w���my���^ǶࠐPwnR��[O���_��PPs�̝s��������9�i1"%1g ��P��m*8�#�a���gyKԇ?�:^��;Ҳ�(�i-�(�pK��z�� ��Ksi̓���C�F>aR�����|�P+�O|ӯ��1 y.����j4�hT*.���{B�# $�><��C7;��~�B6��=<2H$wN�>��#�?���J��5:4��G�E
��C��E�� ��I�����4�R)))EI�{��d����\$D�h���������=��=�ǫ��x|sBj1%��ZhmP�"L�G�)��N��./<$��]{��t��C֡T_�>�B���K��Zt��������YH���:�"=犟5�Nh�Z(�����@�{{G�oߦ�@s�Qf���r	��9�
h�z5C����3 )e󍅭��(���σ����c��4�5���k;��X,�V�M�>EH��m��͹n�&D�����G���q��7�ϥP@��AyO��H�h�9֌l-5�)ր`��}���7�;8��2u��RV٩��KbL�=�)!-=9q�\�����p�~�4����e�|(M�k� �e�\,1�>>���Q,����$3B-��}TY��_\��A���ҕ+�[��-w�غ���H k����6J�4����7#*#ceGM�_o_��kv�Q��5NR�R��=�\��a!UK v�����Q6���� S.����{�I�	;qV�*�����*OD7�SB٣�A�M��M�����V��#��7��s�\�_��p�^5d��X�\�Ƹ66$�)���Q��h���ZB�z���z$���A���QFbSW[��d��IͻZ��ݵ5aaaP8�G��_���S���$�����[?9&B�>�o��=����<==���Qዽ�e�]{�t����������:t��L�u�q���#:�����1'��G��>�}�B�j�n�	��� �=�3R����a ������υ�U�n͹K:��d�y6|�u�h-J��R���xb�sm�,��KW|��%�}�*0p�Y��e����@�r��0J����c��}�s�gg���~/�olz���
{�T1t�E�[+g���C_��L�v�V����w/+�˥�h_��������4J��5��*��������w�ZB�<f��;���X��!mTH�>�^�k.���(��������7�7-w�@5��ǿ���#>Rn@���@�H(gB&��"OV��4@�ic������.;i~AW��º$f�>���A.߾�b�����Z�k����NH�G/�H֌�,.���ArK��ؘ|e����> Q�f���>s�o�(j�C�TyW��s�Ld�:a1�S6���R z��￮m�������^H5�%��B����
z���c-��-'�r7;��G�o�Uv��	7�����*�ں:7�lĿᗝ�*l/�-���)�᝴ް	��˷�2��>�zP�|�� �l�	@y�X��}�Gi��KK���"TU��!m�ޥ�p��4ܡ��m�d�{�Id�����Ş1-�!R��~����$9�}-|�:@���a��c�aM!�s�^*]�Wn��Z�R)�����#@O�L��a)�Ť�qx�_�,Ss�Q�zʅx~��`F�؛�n��=U�?���<��E����o�\����y&��Ũ*�
?.���N���������+Fy*���c�y/�Ȧ��Yq�[[�E��Ѫ�÷����U�I��u��P� ����s����ES�����9U�'�M:��.����٤4�zђ��u[+��G��v��� ���fz�Z ���T��@yK_Ň�4YQ�F���]Z�=Bf���~-��op}x�<ћ)SӘ�rp�A$~��x"T?|��43cFP�W)���X��da���7er33��"dܾ[~�ڽ`�>-����f?R6����L�ES?���ݾP�c�oO�����c�㬻$R�5��ܳ!&$DF�;���B���泞��mmr|��bY�AWFK�*(f
�>��=�ҟ��.,��i�Z��)�A<�\�$�$�+A��~�G�(�DA�4�:�J"��k';�@�0��R��TFF7���$���]�"<GW=��;���2�F%^k�M�̻�#|s�<2�$���oi
y*���'��h�H��yb`4C6����b�H�Nii��@n��ܿfQ���}x�A��F��{Ș���T�}�3'KJJ��~! �M�����]<7�B!ޫh"x�� 
aD\\]����r:�y�������<T��=�n���	�S=�Κ�G&��p9��U�u�#���7�brk�*U�#�%���~���X�������X�[�5���|�ds��n��p���t�xr�?,zZ�۳tYۛ'^�ʠ�:/elf�;�D��R�Xy��aN�&&ӿӦ�r�=c|�gq֍��W��'�z�
�o`��D�x���(��GB��J���8��oR�OI��!�82�2��!�k7<����9ɩ'�	]����Ty��z@}�$}^s��k�y��컦��W9��7 ֢v��=  ��[��J:ߩ4�EɎ�(��ۄ ��]	Cs�R*R�Nf5���0����sp�Ё� +{�-�Ħ:s�θchHVe t[�%�[��}J?}DL� 	Fy�-F��4�$RL-��>*�ы��1q���jtRAq#@����ne	���z�,�Y�BiJU�C���p�����1�v�� ����O�Ɛ��~v�f�L���eh������y����s6�ڟ*3�`h﷥Sg��t=U"�*f�.X|���oF5��h��=+1n�s��*_bx�L�C��"�$�Cx�\�b$8i",�	"sd��l''�9c��ûl�!N\��~Gq������8IZ��~�=�m���%�Ɏ�v��=�VW���W��vV��lXqqw�X��W��>|�G19Y(�]J��ec�r"��KH�W��b�P4{��y�Ч��Q.��T��3
E�,i=��'�� � k�E�(�򬌅�<��lA�*º����)�����Q^��Ł�f��e]YFrĞ�|�)��n�43����#3�����uY���%�Y�
&''��peh�L��F�r��ǐ�Ώ���,.CD\".)s��4�3�U�xe������3��	���'!wh-��Z�+�e�h�.�$�\
�@�īv�&��)axg�4��T����O���q}��q�g{/������3e��>��^;;�tE�̛7®�'C-��1ǋ�$�b/æK�v�hѓH��<� ��:�$s�*E�������'��^F�?�a��:l�ӊ���v��z�#�s��q��R�����ݷ�Rl2�����{�	kB��Pc+�|�T�0DɃ�^	Vlo�������b����7��P�'����k�E;�O��{r�o��4G�Z^PS�ݩ�w��o��:O��5Uoj.544�\���I��l���n��HV?��ə3���"�CG�!"&6v{5��^��M)ᶏ�:h	6y�T�C��͆��B��~{�߮����>��k~s�9����ȧI��5��hWuu�X��߿g�G�[�]Y�.t����M�Q��1r�q/���ĺ���׳F��L,zZh � ����9�a@kԉ�y�睏n�v�EEӻˁ!6�v�Dw��!����,^��_�
"O���:�X�]T$!#3%>�҇���)�cP��.�8D����Fˬ�r� �%ؔ�3�!ӓ��R���Gꅖ�Z�<�<���C��4�R���w�������M���\�m���B�^M��r�q��jN�@�����ͷK|à%��7d"�SX���	�?�`��3r��ǖ6��� c��-1-�	,q�>$�2���;�H� �}U�\>5��P,���pF3f~���	���pUk�� �r�x��p�U�u���G׸yKyK	����?Vy����T#�����8�3���i�9W�T;Kvzgg����$���hŷ�q��?Kcw��.��V��͜�E��.6ʷh�!:��`��M*b̔�P��"��2ҩ��pv���a򡜞^` R����������'�w�^�9O��i8x�7w�T��9��{�/=Z睟Fq���>n�����2���=;���ަ��C��g������L�W��|��������(�&?����ɮۓ��T��4���%��n���8��-����E�Va���?�{b,<R��<�]������&T��� il�Hz����[;:�rtVO/7��?D��L�λ��_�[�5�����sx�>O�P;%��n�����v�(O<)�wN��Y�D�|��T�'
�,T��\�G��&)5]>��A�g4+�%N��S�A�٢]�)�'8���Z�΁������wD9cNV�~] � ﲽQB��qj��y+(����	�:�C����}�� i�gC�K+k.�Zh�I.C�V �o���H#e������888��{��E��/zά㮸H��>J��95uĭ��J6���f"���O�������)�S��-:�B��������lP���q�Jf�Sǵ<�y�����O�Vb��z�Id�b�h�A���|
l�>�MX#ˉl���U�(-�xd��/�=��7�.�Ą"ύ����A4H4s����hí�Hv�j%��7�t�������O��{���5�z����` uδ]��;���;0_���&�g�z-����%~�Y��q%����TĖ�ϻ�f��>y��٠�/���z��}ґ��V;�����r̵�����������Q@@�C�"�y��BUTē���_g̱5CK"i`�44tϟ}о��ۻubL�c�pZ��aO�q�B�E��/o"ۓ��Q�9q�Χ!�V�N꘿!��ʊN/�<
#bI���LN�) t3�.���8��Ku@6�5�#C�u"�=}�/��!Js���S��{@z��y�A�K��a���i⯬�!��H5`5dB�zV	��,�_��	2���</���ےC�=��Dx\���c�9+����˾&��m]]�����ѯx-.v�"^���u��f6
~�N$2~6H���~0I���Z���yņ�?�H-,I}�IIdΞ��Ӧ�bO����<�_�/���� �x�ÙF��V6��I��Gয়:\��G�i����tTU�Q�Sj�.OMj~�Pe$!)�j�VBi#�\��vQ,���\��tsg�fcD���)���>�6�`y	�{��h�LT�[]��Őc�f3*>��δ�(�w=��^J��	�u�މ&�X_����s��ǃe-��ς�cd���TB�l-*>�Դljm�ս.Rv�H0�~�y���!w�X��sN׿iaF�d��
%On�N�x�\e����L��|�KW`�*S�a�l�B�г8���Sǿ��c��5�V�IR/�H=O��3t�Q<�������\Xa�������S�-n��\��B�K��IP��m� �&Щ��n�Ik��*�����fV�J\}�����/ڋ~�+@�7��Z���YO��便�����c��<vuuM,$`�1r���T��O7����q�$]S.�NN/�2s���7dd�A|ԀmwƟ��9�zI
8kA���B \j4���e�y|Ȍ���Zc����+a	�\��}>���~�T�������i�D,1��\4'�B/���}�{�����Y-/���u�H��0�Ú/�n�ꨈ�+Av�T^}���BQ����v7���y�����W[i�RI^�Y�:= 򷕫O�i?�G�5�nʠbxi4� �HIz˿���A^�#/+<L��M,tl'<�4���7�Í�!T�1��'??�MTÆ&�����P������b��CflU}�Վȷ쾡G�}��_�`6��Ў)�m�L��dP�l0�땫�����Ӧ9��`"�;�"�֢O��k
+��j0$�<O"��!��S�޾�s�ϖ̴����7}1�����?��NI�7�<&{��W�Ξ���>���d�tl��\�ׅ.\��?��r��Q�ԉ� uP�~vF���fcN���h�j@ �ܧ���0����؉c��n�~�7@��MJ=��t�9opm:'�yXn��SݹS��z��YGW��:���g\y��;�R����	�D\Kq1.��s�$I���S典jl�����%��0� ���n��R��k�w��m�`U�`s�3�	��~�3��ٯ�x���G/���&����vv�/��z�n�0~���m͈��RH���Ej`h�;���,"����R�.y�;�������5�Ҷ6��C	�4Jհ�{�����$(xk�GH*\�l����ec��W�b�����FZ�Jj���ʚYX8E��>�z��x�-2h&^�8Gb4FP��
����.շ�HQ��l�>���"��x�-��a���?G��k!a��*=,�oo�HM�Eu噒��^s��1w�����Inv�}J��꾪:$Y#_�i��|=r`�.�F���!�h�7.9��1�"�߬
�Q�P"�ҡ�_�UF������XGU��W�����uf�/f��?��[^�PzM�H!��އ�O[��Q�go��x�Q��2�T��t��鯤[,�r�$�>,"7���i�,ˁ��(oﯸ�_`�C^�s��WINՌ����#::4a��P���������rW��k�k=%W�qd�����\����WMmC�"r�����:�v����^���2�Ts����GAlQE�k���y�V���3�I���B���3kkt~�Y|�γ�z�1S�Oo��sʾ Zg�C��*��d��������-���M�E�*M���
�_(i�1�W�eukF���}���UK_��y�x�t�)=ނ	9�����e�0�����s#5oب4rl�]�F��p��eo�Y�]�v�%t{��j]�������l`Z.�o���-��7YW�)u�L���\������f������(hPd���Eů�P�8��Z�k��A+�ޞ�[X6s��xK`�Vvt�u�[iX=���;�]��0�u�p�Je�5�R�`�b����oC�cD=6���y��2���;���=��P�u�,7EY��~��x�����U>�o���/�5W�#�7*�k���������U	�awo�T�q�=D�+��7Ǘ�s���=y�|h�ݳ�-ON��)+-��̌�+��;��=bb.t'��ݖ��ܼZ�zQah��E�W�TJк2������Ӡ�@��K��T���ہ����:�={
�Y��17E,�xb��0U��lxg;Ǣ�Gs��QXC�3�{5Q�9�G*+{�H�M����ÖG�G�(���p���
"}�;�ǅ{{�tŞ���c�
����>��9�O����>�^K�+�����E�����nHL�`x@�&ҽ�`mxТ�����K���-�t~˔z��ݨ�w��3�W��]>��y;nu���e^:w����ΉrEZ�u��K�<�9�>	P[��ޛ����|�'ǈ�(��lq�q�2�����O� %>*'V����r�E?��Zv�
A�񴂲OȨ���u�]�7��S��햮�]��]Ѱ9�!D)�y�i#uL�4�C����|o��	�����p��W��ǎ݇G6�Gf��<4�U=�r�)��+&"��O����4;�l�H�D���BĴ���ciW�i���׉
�x����������g�w��ߟ|���E8�y�*��e��b��mQ|���nT�2u�/N-�8��DV/e��AV'���"�\}(He?�0?��U/��h��{{{!���*�_�h��~��? �X�s�����4���!W�����K,��o���dc4����]�o�s��l����mFDs��+����{�p����e�
�������FZ�x�>Ř��V��$Z���0I���Hѕtr��o�-D캦�<O� Wf,<{�l�:���KQ�2����kT:�ݳ�yx;��q���<���v��5�ޗ���=6C9�C��"o�p�Ցa����i/�}��Ἳ��NfO��P�`Zj�@��S��� l��3ٓ�|�i)t�������� Dy$�����|�)������2��	.mB��u���ۙ)t�#=����O�<F��S�64�Vz�+�/]�r�P���pJA���&Z7��G�x\����H��2~��IX�&��Gם�TѧhTI����KR�F$�n{�ܫ��&8h���j��I��H�C҈��a�P����bKs���~���F?ۑ^5���*V��uI�+r���2�K�����n�R���w5}1�O���˛g�a���/o�4z��5H9o�>~=�&���,��Px��� o��2�E�Q��G�nRo�qxyyk�X��p��EZ\�wɊg4�OM�/̎:]�����Jn+މ:��������w�Iꖁ�e�
�_�4�^o�X��n�
����`m����(��2�H&�p/얻��ȺϾܼ'0R W��x�/eV���&������?�f=��۷��aD�VUE(L5������U%�]�+8=9IDI�D<�̂vE	՟3T��)Ar�W�1x�M:z��k��M���1=n��ѱ���|P7+W��ip�����o�Uo~r/�ū"ss���i������w����_�V��m8�-,Ш��L����뚠���'&��+���yΫ��@mz�z���Ąb��ڛ����{�{�����|s�5L^~L�� NZ�f�a��]i�^J�I6NN.��nd(������|d���:� @��o��ze�+��
@Q�������:��!A�����/\�;�M#��I )Ҍ�)E��7�cE��+;��Q'�F��_�9"�m�����J� _D����u�N�E���*?j�����;�W���qJL���♖���ݠ�Τʨ�9`�����tQT������~=l���)�+^0(�&�g�:������̏��e�Q�i��c ��Ҙ�G��� 5�mn9��FY99Qx�~������:��ӛx���xc�֖�Q�Y�B�?��#KKO����)���u���m(�#�R��}/}	ZEW0`yZj��īu�3��6��ܱ�u{?��!5|;�n6x�����vM�v��5������=ы�?.rTs�$�W�c_Ot����)��il���T���]]�^ƾ��"�;�w� ���nD����ؕ�Ţ�kj�aD2K��e�p�U��i;��:���gM���Ź$-��$�Jku�⩺^��3�$1��Bl�?��z���d*$$��^��(���hۢX�*� 6�;g@���s�u-�_�V�2R�Rg|��W����߳MB��I��I��S��ȝ;��)�ߊ�v�L�)@w���E1�wm�I�b¸��͚fW+�t���
Q�Ǐ����)���O$�4��#9�3d���Kg�#z��
{5����G����DPQ�Sh�0�	#��ߵʄ����%�j�D� ���2����s�N�~�`0����$}�.]���U��z���t�[�9m�\$��p�����L,�?UԿ���X�ۂz�;_{U�
�GR��`�k�.{���]q[�!૷���}ۋI��J�N�Y�S!d��v*111��@�%�w��}ԥK���w��R��� f���W�kk�HP[�{��rpU~�����D�����'we�;�z�4�N��F ��g��$�D�@�-�ȁF�*���+�6"W��s�ĄM@t{n\�_|N[�+/.����Dn��H�%��Fw������m�?�ϑ
!n �z_���fN����e|�E��&��#��X�(ص
h�aV����Ǧ\��rb8����8���ъ����0OS���&��!����ܡ���`҇�j/J�؆��>7+I�:�����ss�Oό$ugSFK[���u<H�M����Ύ9-�CJ}�m,Q�,ӡ=��u�+�%D��p��(�_��k�T#w�c��?�b�� �i�3֯������c���y��꾖�>/+��o!������S;;�

�E4�\�|�"s��<�c���%�ʅ��J�����:�/����L?WOb2�m�3ر�x���~�mK'�B.�W�������r^[���o�����D���XkÎ�i��ץ;>MOKKc��3-��Q�m�ec���k�����y�k��F7ve��A5Ci�&X%�k-u��H��.iEE���N6�8�UK@��ܰ}m�{$��I~��󼻅��1ᔦ�N��G���Z
�8�<N���P1���/�Z[#.��	��TXݞ\ߙ\��>�V�ks��)����Wo`���J���Dk[ݿs�_^��u��l;I�fH�~u�~����P��}�]���.J���g�J��� ϞR}���'��\a��)�-�<��Oy]��/F|�ȝu�JH����/���tt}79@���Ni��`(;A�;�����V���|����"�O�i?[&�raF�@L$�W��!����h�-�?b_=�q�exD��ۂ���(�F��]�M�[�IE%+M�ڙ��3ݢx���X���\<�y��<�FĂ����W���y�Ju4��}E�_�9��i�c�ַ}�"��%�,�H���ʝ��e�̹�|�c��^�Z���Ž�IT�\;2E����w�D��ӳ��"�X����!
�	W����T�B�`@0�~J�YG� t���Q{~
'.�&Ǚ��r��w]]]��7�s����_"]�z	/zץ�$[0V��9؉�L��n�~��ѣwp���]Ԭ.�}��=�]T �$$>�\������*�|>�#��`�x���)��ڱ��ص��BLV�����d]i������Ab��臃��XIM� ��h������3֞�gdM/]�ߗ���С4�vF6������q\V��mU{�'��������I�'��t��3�7�cPZ؉0��N�c��#e�&Dp\]/h����� ��5��:�g~^�%�m�N���'��R cᑟ���m\��A��,����+��Ñ[$��CDi,�ߥ9���x7<�	�`z�+(����_��,ͧY�t��������w��.Pdɲ�lr�NM�$��pwo0��u��{��A�&���Ib�-��AY�-�	�p���v�~�f���Jm|���xE�C�3����g@t'#H����Av�8�At�.�7u����<Q����^T#t�Xms���0��u����u���v����*nv�&:%�raEZ���XX"��=�42��8z]A�rԳ��^��Z�gh�[|�.p��_��֍̒���y��#�!�����.o{�n����S�Jr�1�<8hFl-0'ӻ+%!&�}��e�g���:�$ȩ��ܾbm8Ψ�j�h��r�EE#����=��"���,"&v�� ���O��{=A�R�ib?��_�H��YA�����{�1v;o�G�Ȇ���I��e������f�{y��;�op�f���2���� �B6�^�s�~ّ��7��<e�����)-�	9���W�V�TBT�p�2���M��%�����nu�x��}@hη���>�����rn�}C�2xl�(���P���?t�r���pM�I��a0�	�)�w~���ș�r*��I	�+�RS.��G�%�Ƚ��c����_�x`�X��;��4䮫<mW<�5�[|�h��F:Eѝ������/j��
[��O,w��H	��*%vv��6j�s�S{uC؆�Y�<S�ck��f�y�~�5|���Φ�<��^�3S��>xŮ\�-/���+�Qr6��/\���a����`8vM6�siI�@�k�M:����&�鰥�%?�p������8�[qY��r[�Vg��x��'�U��ʫ����m�;�-6-� OZ9��:D!�
\o�ȢӶF���3�;/��g�J��Cdx^�8J���"WzO�UfP�m^C����[[��(�5����s�d"��G5� %��(��R|���ff�k ��j���<�H�u�xOvw��a4�X(�GT��_@ɛ7C�ẂIo�֩��J{�^g=l2Ev}�Rz��t��)~~T�P���t��]̌	߉�U��"O�W�l�;(�|��WO/(�u5�s���s2�P�V2�7e1�X��1�{�+��%<2��!]<7.���fy�	&���QdG�h����˛�"�����s�\�	�����;`j�N*0�ȃ׸t�^�ڎG�1#�/�=�+�cs!(rS���3����yDY��ڬ�"8&������S�j�Ґ<�;<Lb,�R�cTYZ
D�⇶6+3s���wl�pT�ֳw���q,��IVK V��.�ۻ���18;�?\j-���m�dvfIɩ��$ǈ��rs}HYF(8R��1(w�'*1!b�NW�����<��-!���}�(�FӋ��!����"B�g�H6��1����=�0(�XN9��9GxԐ���nU�Rd�ϩ���J���(,��b	]�CFA�)���� �m�����!"|�J���I?�A��0�	�H4o��-=r��Ŀ5GF���!F&
�"�範w�x�P����Ҿ��\�|>�Pط_�fz�7��5ց��[����%N{�'�u��}�x՘�c�z�S�]0�{��G�TBQ����ɭ>d��t�1̾Ѻ�a��)�@YTdi5�Tڵ��~|"��0ӶL"k��Tǵں:e�$?����O ,����zx,����RBe'�HI��PJv�ΖU��3��
!{e\��I2.�2B�&�����|����qw��q����|�q�gˁ�\s���3ˮ"��ñ�/�w\�WN=4�[�w���R<��'�Ali�-q��4L����3����|6����w@TN���9?��� ܌����y0>dN�����F��&���FZR�j��j�`YV�f��;��F�N#K���f͆ƞ�ж���r|��m��^��_��2X��C��/,�X��z.���=q�k���^��� �voHepӷ��3�x�ȃ�PLg ��Q,�P���Ґ�vp�L,IbO��~qdL,�KS��&�J��}��e�A٣:LE^���9�M Q_����m��
5�?x��="�#d��BYp=�+Z�`4���PUZ���v�A4���!�Ǉ��>��cR�jV�{2ȫz���?�T�K�d󹗭2w��i�m.���z>{���K�P#�=4o���c��?~-`��y▴x��%-���������U�pk׺QP���b\�4�4�̓�At��nq�$�>�͕�f �i��&�`j������!b|@��N��F h!�$�.U^^�`���[C���!k8�l���%'�O��[�΋a�m���m���Ӿ"oem����76���W�F#x�F\=_�����w����t���;w�u&��/���v�K�w[T��e31E���E���j�|.*J���-J_�y��I��T�)5������EZUu�O-id[_�j)�U�3�N|}|�l�o����qV�:55uNSK��er+s
��j:5^w����ъ�H(�;����� ���Z�K���|�P-0=��HNª�ȍu�z���5��G˩Y�þ�ö���>�y��A�UY�����J,L��!R���E�ww)���l�������MK%u�F�!򞨻i�����JDee����ʜ��`�N{[1H�'���������n�5��[��0�ڃ4��Kn���=y�����6��>�	!!�@u�����i�����t/�3o�s�}�8Y��<{�J(�%��Ը�*7Z��[]9���\��~	D199�S��	Q�y���R��v!S��U*�9�
�ZR|�'Z�WV��T5�3Bڅ�b(�op�BCK+��r�P�ZUٝ�D"QRZ���W܈JW�1��rN�QdM�!��pCs�-�"�����$���dX��"TZ����B����������K-��e�@��2U�8�REȗ�j���q�w��ՠx�&�@�Խ���%��W>��^���.��q�W"�����S-ky))uuyEEC//�荏��ے��<uby��+�HZ� ���8�|�SP�0��~94T��f��=�<O��{�m����	Uh��J�G�Q2��)(��3Y�er~%�ć̜�;��"�Y���:F�~��[.N�W~���r�nٶ$d����pF������Y~&|����|>>�s7�̧�q�*.��$	�K0특gm���u9���?M;d(�6�u
0_C��eSE����}6�o7얦L�
�x��iS��
��@SWiJ�����\v��^��sp<�N���U���j�?�P~��ia��+O��-��25�����&�yq�U��\&�B	S<m��^����[6�B(MN*m���]8����F�tӃ�����K2�$��������c�g�$^��*�ѧ� �xmz���̪)���sN����ww�L��]��DDD�5�\WTf�F����cU��p);��$�p@p�����N�y��h!a��ؘ�	��VWC��h�=���h /��.p���1��:���
��^��ӎ�vT����4�?ͥK6ږ4w}�AF(9ٞ#���'���������k<"���J��쑗�ކ��a�ݙ�;�� ������S���l�va����s���_��U�kb��˵M���|��t�+'v=̵-���8�M�\�)���I;'�o��>-�a�J{eZ�����)i�2'��}d%���}����I��Hq�X�ֳw@w�.M��$s�t��Ȋ����QQ��$'add�g&'���O�Mk�f�T���{YR�W�5wF�-@���TqqqāV�7T+�I�_o�y G봺#������$��'�sJ�T��a�F��-P�w#GG|4��>)�Is��^�11~�����1ί2�)\���ʊ�Ҥ��?���V6n:��(7���<dg/�{���'o�%��5�!��Tʻ|Zr�6��앹>�� .	��+���L�}��z���7X<l��8�%%B ]V������~%�lX��C����Ńmg7~�,���kHE_�xꜝ:p�}_�uO�C���$��_"{5��	1����ȷ|o�^ ����"����T����Ez		��R��|�����^��an�]:)�H���l�3r�we�{m�����Q�VB����nq��A��m*���|/{zh�;��j���C4���'^^'pUL*f��nz�9F����Ĭ3ŝЖɦ�=����555� r&%��.�J{��+�Tc3t\�*�ML�,jci��,�c�{�3�\�o��ɮ�q}�fWÌ�����g�e$㘽F�=���va �w+�����ݼ���l�Z�т��?�W'�[��8�WT1�!�Ȱ����`��d�9����nk�׊���C{���OC��`���L��ߐϒI1ʂ���Rk풙�N����v��z�e��zz4�y�苈����~W++�Ț�Kڲ<�	�]��Y$���5
.ęV���*8�3�߱lu�k&?-idH�'Z�ᄺ�5�����;����ыp�"΂��}vj�7�ODw����~���iE�lZ^I�	���3)K��ic'�5mkI.��ܶ=�)�=�g"���v}=���я>�vN��K߀͵4����B#L*,=�B��R&��R���ǋ�~���Y�_��,���[W�h�u^��Cd����0�QX	P�.Jq�?��F�%����t\�����������L`�]f-��T��l4Eh+���)��cS��Nlmo���|	i�P0���܌���Z�C�༕�O���wR��`���X"�e5)f�e�_ߚ�_��M�	)+;Gt�Ѹ�6g���X��pUƫ7������eh�/�dO@Q4�$�U�@`,�0�g�{�Ė�(u��߿V��b�DZq<Ԉ*p��Ar���8E�����Ld���g|��տ�o:L�SR�R�?9mh����y��ѳ4�ŵ
�X��5�����������É���(���I9���c�gY��}�*��*B:�8��\Ƨ���H�F���!i�̺�Rb���P�|`�a9�
��DK�2�簢��%K4%*��A	��L&��hå􋗵T���6��qC�� � ,�L�
��J������+�}|RL�1���R�������� �k&���Ȉ���mP�ᛢ�F�*�h� 	�~G���5<�o�zƓyh*2���+n6%�(�v��Os"�:����{ɼ=���k����&����wn�@�O�E@�����3F�vF~$Qz��Y�C��u���4a0�_>q$E�E��##�^bʿ[�fp��j���uo9�a�����~*yy��<69�V���!�m�\��ː�N�r��)�cp�
�2硺���a�H􋱅�0�b	��3Ǉ�,�c�ojQ�_a���UP`Y�8������$f?}ͣ�ܿo��[�%����%�>3c^k쟻�
$�0a5q���e��.i�N�f�Ezp�B�|��	�]r�O�=:�$?57S2E/C�rq�B{>G�B�����e wIEE@]�a4�rU����kK�m|��DғQ���-��U�B���>�h��K�։�E��P��''f�IO��FB8%дϘ����Al�M8%��v��X�3��׃�������-���*�gs��/��%��5LL���p��p��T$���ߗQYdi2��:4tb�2눣�H=$��MW"0�����i5�X�,��ȶ�:��M�_J
���R櫙6�5#o��K뱄w:���G�������)��኏��yn}�k-ųW��3���W{�Ï6_K� |�����Y4&ni:<�,�"ě�5���j�@9U�g�O�S��S� �ύ��E�����Jd]�G��ѝ���>��k �fg�(�Wf����;�YJ��U���1S�Ǝ�b}��)�����)���]��X�P�;��T��B<���Tʏ��������6q� ��q_�3�'w����"���������6��"o��V�3���O������s���ع��𞖍�9M�<a�������&�"	�-���|��������H3�G2.����-��<�И񆔪�)�����-�m���x���y�mN$�gς:%�e��p�/Ҝ�Rcޫ�b��u:&������¸�ۧ
پ#�b�l��--�	<D6x��.E^(((�Pp�pc}��J���o����L�N~_����e�<�?0���;#�Z7OO�p#F��8'�$>�������M��A-~���uH����{�Pc����.&PE��9�����`ck+�:,���hd�YpQ�A��5p����&#M�������V!e_���YV����r�C		:�p��d���K i�093OS[�y�����B�̵=�Ĝ+�����*~6Zŋ����W�/e��y���)��t¥�qN�j!H�"|��r�DW�E�Eed�t)��4��I�8S$RY�M�-��&��B#�Y���:n�I�����;YP{1��zD+?���%F�9�pڱ�i"�<���@RjT gW�~��c:�{V�%��?�2v�U�+wŘmf��o������n�{,K�WW�<"C��ea�gf]��07/��8��j� p�&p��vYv�B�z�"��ee����f)U��^�8+�}�`}}����`}��S���n�"&Z%�#������rװ��J��݈{M�]�����}9�ސ'��E�7[׏P/Wʞ����9h�d����2uOh���,שHk''Wfe��rM�GGmm/lz��_�=�{�-i�TR�i"At;3e�EEnU����_5�KQ���w�;��_J�zQפ��MO
C,�k�Ȃ<���m��_&+r7<�Yc���^~':8/�M� A�o߹���� ��UfrR���d�$��q�l`��HZv��U�Z�8FO�hp$��u�c0�պ6ض�翋���"�F�̲R|���Fl������!�pr�c�:���5�Wȉ�����*�yuD��_��1GV�tum���j^��X����O�gCv���kR�lF�^<{��(�s� ���������zv��6)�� ;��6p��xa����l�O^JJJ�V��D�a���;���`�y.�������i�Mtܫ��Nf�������)>�vj�܊G=�� )0Αw��UU��&&�ߌTES)T��+!�C�����*-��jT��#�<L�*���)�Hez��� �<å���p�������N�R�g�E6�W�<HrrǟXXk �X*+�f���Rm���R���u/�2��tI��+�=�� �6����|a�&�71�+�!��KM?�����=��xz�u6���'1����tƏ׋�/Ʌn�Fp�.F�������C�D���%%ꁕ�e���ihh^��o�Պ{(|������ERXz&y�W_�"�����������%)�x9��Kr�QPϨ�i�3�扅�Ɋ�����5�ɯ�(��~��$INGNp^H��#&!���}��i6����DF..���g�(��S<'~wZ�����<���7O����4���+,�������T���3�&t@kt��.����1��M�M�N{����7�$δ�J�N�x��85?�.А��SKs�_����"��of��QSS��HX3k!��+$h���4�_o�ޏk<����<�3���<�	�R���!F^^�ف�4*h���m
��:�.�DHJ��%$������?Ń�D �c�^YAe�̵��&�4���r���5�E!Z�m��)�e����n���aLk����Y��[�3��ӧK(=6K�������kP�/����L~R���V�&���-�sr�*�0�k��t��N���(D]o��P&򛚺
z��I	^��r>��I�`3~�C�c0Nը���*��f�+}/�\�
��Y쑻���HAZ�3����j�BӃ3��(X�+<�gi!�z��Ċl�Q���u�ѥa����Su�JO��+J�#��m�r�8��j���� ґ]�Z��R�����������'�x#�]^�+��69>0 �IOjlmݲ%a���(�96&�cn�;M1�,{f++�%'���B���:_K�p^SV�3H/|�u|���xŞ�N��V�y��M���[L�L��Q�y4�EE���s���cb��y�6:�;�����}|��?p0s����X�&�J����=�lj�N�۷�9[�~�
而,���L�0��[�Bݼ>fO�&�<��J�V.���Y>�n��	/�=�r�)s���:�Oc#��oss<з��6Ų�N���fv����kA|��ڨ�ff����­������C��xD���M��jt���8_���P��nz )���?��w�ɓ:'ffhw�OQ"��>������,H��3���'�,P���,�g�cۦ>���=T�rt0�{���,@���iʐPă�\�JII���M���"���E}$�dʧT7��"���b�s��|E��g��D�C�k$n�9���a��S˘&�����)�7٤�Y����{{�)\��o%Ì���R���=ill�����\��6	�C��	�q�rDF2�-(%m��[Ȁb�=ST\�Z~�n��Y�%!a(�Zy�B���R����;	u6z��n��@��X9$�n2�����^�z�(R��3�*mx��(��\��?ҙ�oXm#8c�Z�l*�	Z9���f/�H�B߇���q��ȭ �����L��
B�R �J�L��ՠ2��ui����ћ��<���������z�:��I���٨#-�t�0��{-vB��/�B_�v\��'o�_���O������F�*�P��%�v�N_	D�� *�l���*�O���/����9�5�4Zt��;�{�VR�,��lZ\�`x��x�FQ���s��*�r�O��t\�5)!Ư�(������<�:�p*����Uف��?t(z�[P��.�O�-���R��`�vBa$n���6͸��v���+/͌������[g�Lx	>��y��FA�����k�����rvKNⶕ�������zI�&AV#w�S�����CK�s��H��",/Y�@#�a���ڃ�s�� ,�Z@X0��>Y ���B�)1Y��"V�;���w K%3�Og����w�_��q7�; =H����1�/8�wY��`z�E��|�J�t��8�=����n�11UG��݇ ��=�����~�0߆c��#�m��uL�z\�q�(��"�P� �olj��0��+)+�J%32��T��(����-V�`j�[卋=��4�.5�Ԥ�tC�Vh�TU݀�{#�|�uйL��e��Op���E��B�c�d��^Bn=�*�`@�����g|��'*6m깭�����> 9Mg"�_@%ي�d`��`�F���3�?������IW��Hj=z҂�D�p!K���
D�\."g��j`@��ޗov�f��~�>��T���%��JRg�.�U*��͕K(�?f�9�{b��@z06����M�.��K��O�Ѕ^E·P��A�AZ��4���8w.fe�_e�A�J� 2��Йc�7N]�y�� ���U�<i���nbHP���%��|��C�؊��y�!	�_�F�pM�i�aŭ�w�^(��#�?ۆf�s	$�6�'��A�,��/��-�Q�p�9-(8� #U�e�������oz��=�f��7a�_K_������?QXߐqcm�^M���Io�Z�p/��$��]R�� xV���w����>c�6�AM�5�bi���FE��40��Zx�	).�|0����ܜ:�o�^�_j�=����c������׌�����9
�x�~�
K��{11�̔����g"M���(���Ln�9�Mc�~Kg�<&��Wc����������{)��B����OMx�e-LpuC�8 H�:e}9�|��Y��}� ��!����W��}��P���s�"��+�U�E���
.�K��)����_�6,Z8[����_���U �&��[�5���GVS�o5���/��n���x)���;'g˴C��������o�QxX�e���������,�����b� g^^��	`�I%�~������,�_��sml�d�eO�cض�\n����w!]ݩ.D�~��I�q�:�L4�^��n���H&]^'Z5I�1?R ;���4 ױo��֊�.'Ϭ���G�]���b�{����ͤ[C���n�B>Ͱ��r'�z���G�H0��&+�΢�x���٨_�eC޾=�I�.�磕��]k��|����ܵ���f�-`+߱�X�_++����Ty�M����6ge��lnz0 ���b��Â��=FE!'"��ڤ���<����TŃiPc�,��롕�pʑC�����!3
Z	6��^��Ky���&d�O[G\�s:^{N��a�lY��@�^�"+?Y�*�F�]SF��o��Uy�(�Q�H���o������^M�n�S2,�����w�l�9�n�k���ײ��w�";��ؤ�B���]��5	|Ԋ�G�}���e��.CV!�%�x��#�<���%���b�nP*�d$-;��c�����bg� ��׷�������C������:cp�z�<�����Fl�C������!,*�C�҂�	B;��`��)+�I�_�g<�z�_W58��Ç�k���w��jZ�n氞���<j�����OP�e����E�����h��p��m�$�H��-1~�������n����Ai�r����E��.��ۯ���sd�m���c���������H@^�`�MP���W3�K�:Ս\�S$�S��SPxc��h�
0P�Q�c��;�!òq�ab ���	��h�ar�������>��b�:#)a��p�c����e�,�ۮ�����''��E�(��;&���#�z��:�d%X�
����8�٧�'9ȉ���/Ȟb��]Uf��qQ�SyCHpT���
�Wk�G��u��ō+�!��u�Qnb�/p���#�A{��4���)�������<99��О�(D�-�s,�FR���+�x�����>�A<w�Aĝ]�,+��q&�2(�X�6��-��.^��x���:^43��%ӯ�]��:3C�l\��g��E�[��N�Җ�9;��)�����ÇLADp�mN�e�����%(�y۸cH0,V�h���M[n�բv�a{+��g{���שiii�"r�Oq��_�@���|hll3?�؈���f�����ψ�l9�F��������������/�yT;�t��EE,�����O�-�B^J�Q.> ������gx�3�J�����}����
��.Xw4fiB�bJih=��z�2���h�O���nBa��o4��?�a��Ɏ9�r/�{���/���z�!߀KKE��v��/���ǧ�	�RHT�iƅɃ��wf�Z{��ub]���xO��QZ�Hx���z��m���5���
��vřI��˽σə.R}J�oB�"�O�59����f���x�Y��*�1]�r�HBB��K���*�b}��i��i]e�jӨw�Q�K�^��O#s��w���U�:��yǆFqr���(�G��%��lB����hV'�$j�0!A+<�qUkѬ����嫸���Ĕ�����f����JW��򔒞2,u|||�>}�[���,]N߄�>����d(ѓq�7b��}}=<��95����~���ͽ�Fu�d��ޭ�t{����G_�-<n���̲�?��8�חUe�m:���XUUPX�I�{be$,<���7�3�x7�`�G�2�_�\���B0>
�C���$
%
W|Դ�q|t���VA^���#'�ؿi0��CXD�ҎM����^[�M}�e9mtd���Zr׫�~��[��ܹCKC��{t��UX��ܯ_�Ϟ]4-��&Z|ŀ�$��������@.��4���]�|y�,�ԤG=wk��*>��Ϡc�$--o
���*�^?y��cs����nAX觭�[�����Og��w�ccMk�<g�+��8���XZO�Pf7�F�P�K��4_�i�/ڞF����0��lȷק	��989y�\�$��Z�֭2ڋ�M󲲮Z��pRX�qg���n��[2�������ٳ�j��h5���x�吿677���,�udb����j>�� �7;�Q��N��p��o o�jaaa���IS��6>A�\��H�������HZF⦲_B�:*��N`������)mos�H_��:;����/��1��@����� 2{��˃����.v���I����D����d̠1�Ztt��<�4�	���������)#P�%��
:�J� �BCm.�='�Vx8:�7������ѨD��!n�;KLOkkM���򴆆���\o�e����u_]Aޥ	�0_X��ţ�>S��3M�0��.������P�������z۾V��(��J�O(�D����{�g�x4s�s��b-��g�߳�$zAp��qB����=j{�>�����L��D-��jt��pr��-~�x�r!�38������������Jm�_�n�*�ȘL\�7M�ѯ�(������m�<�e%��0A�fMNR��E�KaW�n���>\���_�H��L�:�B�s(��Pn�Z�I���tQ+��M��柩_�Z�M��t�k����on~aUWi��:kni�*-D"G ʐc�;�ijJ��ۣm�tG����prv9�D8�������?��>EH��V�F��2K���*�f�^ΨsO�wNI�d��J�u��Z|<�;����)hp3�[P���ټ�[衡�	b�=���h�O��iR�^�=�
��	v+mMty�w����ei���g�f����bi����z��oB3`>n�����`�%6�ʍ���@0��d���P>�C�ml���6Qh����v��-�҂�������[)ii7�;f�Gl������_5Sq��m�]�{���%��ޛu�==ʘ�iY�D-	&n�Z넆���?��-��p_������P�[y:
F6L{�*O���sh��`ajǽ�L�v�P>%%E�� �����^����d�~��O+g�����8�郛/�'J0e��݅�?��ƣ;�~7�1�+���}Q�=�C��jt|��k�{�������3с_�<�����͵���'%��[�m3��y�oݔd�ʏh����G*(�ڑ-+s�c��?��t=,��g�:��A�B��ɚ ������^��:�P[��z���Z�v�+;55W�����c&n�LQ�� J��Л���3�$2����Պ�1X,�Ma���W5M˴@���@�6��~*��ө�h�x���D��bʪ�KR�Y���z'��	H��s�M6^����֖��\!{Am|L����������O�蒐�X����_��o���D�gQj�j�� N��M�[�S�c�8�`|��ring��?��ݿ���L5� �53{���M�a���k[_5r|9BQ��E�X9tq񣃃����.Rny��c\�]7�N�Q�gR[�yW�lY�������#P���ng��\���v>�)����+U�f��
Ϟ%d�8�f����޾=0?�����'Կj�LUG�u�������������-�9�c��}$���O��.�v{�!�K��/loG�G�c���
��+�-]\[Z��sPٔ74�ttt0�L���+�ݏ���?^u�hnP�T�,�����B:!�j��R��������
妧�� �]3rMR��|b��[S�a^K�kk�o��&-�������4mu/��SM��u�
e�{�Y�\�A�;�GE"ˬ��VE���Tء�.����< �,a�蛿���7sww>7�����:��|�}t􎶦�0o�ewwwEC��z'B���\�^.I!i��[d�N|��ޞܮWj�7�,Ĩ�9@�����^�6��ֽ��<t[����p�*u���[Y8����_��>7q�"�ry\��1��=F�<���O�b0��yk�g�t����*J��ܤ������>Yl�v�7Gu�����r�1�CV��1˞$���_�W&�3��w�����.]Rzwʧ�����*��Ν�b�s|�Ƿ��L�=9]otO�����?%J;�x4<�ZpY�Ҝ����uGh�ڏ�o��ߛ�
��e���ki�g����8��N�=޹�QZ^���:��~�]/����u��FHHI͝�����@�۾4+��誷����j
G|9�>��t��x�#
�4��d#�9�V���ް;���:�34�xL�6�o``	��U���|�<����f~U�#�Z�̯!chǅ��������݇U��N���e���l�pq�tT 	��j��WA�m.��tu��n~#�l����]����30�|1�N�9��a/`�@�A�g���ٹu���k��;;9��֮��>B�{�vk�t��M���P�S�9�T����eQ�:>O�{ob�UD/�蘒��6�j4+��L����/-+�=3�;h}O8ݛ&0ci�&[�~~nN�w-�	ZYT� ��v]����*D�<K������#�<�JC�mv��ӲoO���z9y���=��oz��-�����mm-}}#�n����R��޿%�Փ�Eu�w\0Ԏ՝b��v�h��f����W�����e,��~�>7��d5�L��8�#p ��D��N��~c��v�����>>`
E`Y��� &��E�UU�vv�C2��H:J��6�+�*�Ch���:�����EE6�</e���h�e��:���������w�3��i_��˙zv�p4�o���v����o~��d��!ꕝ}M+N��륿<�������<@�aw7ak�e�'���X�i.��J�d�'��}��T�Yj�����.k�YC[��z��_<�� ���xl�4��II���ISB�,>z$}���Tέ�'��^Pp
�H�>y9���ޜe�c���]u�dT-*�urO�LOgsrq�(?�/���f����Y"ş߿���p���tvv������x�V��/^������8[.;�![�>Ꚃ���v��"�[.�����\7���̀��uO��2""��-ncG6b���C���,�b��� ½�ի�����F.��B[u�<c�lml�XG����`J�_��I�2�!����݆��[$[��-���w����f�W���[����/���{���D@P���4��~Q]�Ս�'tttFۜ(�|		����uH�FD��9�O�������*��>3��c��oΤ�{�)�q���Tv�KK� m�F��D��2F6�^�g#g��<�=�Q`�*}N0����ښ����z�O�}S��/�VP�od�آd��ַu�{��z�mQ�6�B���Z~2��QM�; X����e?8��zz{u676����M��:��!V�����6 ���?���`�L���W2+�Kl�\l\t[�����`c-��~~Ǩ$�u�A#C�̎W�Y�����nL�j){��&x
���;����E.�mP�k1z�b���4�lԡir�U1cg^�	�l�6s�����������z�uʔ���ط��ֽv�f�I�n߮A�ʋ��z733�?��=�s�{���@
��� ��)����b�HW5g/r|m��t���O����:Eʔ�8���*|W�6HDŞ��������?}q9���&*���C�c}�%�ݷ�&bZ6���s����#����s�0ߜo:wLT����Y�^���2ۘ�2+Pc3�[�)c�}S���l|R�[y>������N�
����m��v����:5࠻���l�N
Ed!k)9�Bv>>E�����ʷ������z�t1������(�!Dun��fB_�w������b�R��ۗ扻���W_�<��N(�յ�?4��=G�V)�M����7'"b��L�3���|*�y{�u�,-E��n-�p��X�������:e����ߝ�FGF�4ٽ�|��^TП�Eu}؊�M���Q���iW�ieH3Z�����Cչ�i�c<�Nnb4??�Az[ |��M~@	� �[������ŧC[3��-χ��G��1::���j�V����nj*k���5�0��11�4GD�]��G��Ć"�Y�%h;��{]}31+����?��������4�i�Bh닻>��nm݋9���ɛ�ϩ�[��f��#�ml��lwhk�\�Q��d��h��Лԡ޻��"oІ�J�{���,������9y{�_����,�l�:��8Hp?��^oqii�1��b`45��@?�S��}�^���	/j��6��p2�����M�+���BU��Y���«S0�;���Hl�1O�Y͵&�Cu�$���
��ؤk����Z�qi;������|h�
7�V
�Ā%@|8ڪ�P`Ѱ�}�ַ�>[�:g��}����ʬuz�6Om����3���K�D���n���N�KIK=}6?d?}svvU���l5�`�I3�>�
�ʚ���/���:,�>�1�t�����B�:�pkfx�=x��iu#�nm���:^��pB�u�0�hbR������sxk��ϝP�B�����υt=S�8�߆�W�WG���Ū������Δ̞|%��J"�T����x���v����.ӭ�QA���[�@ ��c�w_D􍜤��{`��xs?"��k8���\���d�a|�5���s���X��  ��,O�!~��G��M�d=Ī���`S����}�R�m�,Fn�g��x9���SO�)��f>�t��4�ql]�kae����s&�J��0����
Ň7�{�5�7RM���.JK���v?7z%A[Q"b�=�$SU�o��K�?�r�l{���.��H�/���N*���W�F���x?�8#*���8F�&.nl`E�y���뷧��{���Ò��������G�0�-,`�MdJ�i��Qzw�A��aPH�����K�>�/_jI��ha�ﲮf�>���33#�}fB��*��W�÷�o������q�	���;�f�>.��M).���Ǝ�x��0 ����j��a�&�|Mv���>��*��OPK=����c�ӂ~%TV
����G̗��=*�L��Tp�CX���9�ow��O�[��ȚJ�	��z9D]~>pr�����fJL�@&_���1��P�{^�q�(��w_O�J���_�<����&�sa|yj�0�W�Q��a�ٚ����J�?�@�WkiG^r��VXK�ﻶp�h���1��UP��]�S�o<�0l��<�:t,+`S��׍r��Y��`Oԏ��d�6�$�!��sX��iqp5o��Ȑ�]j�v�dis�$`�K�4�t����eͼ�M�qw��侙uo���-bճg��^������p�I"�90H��Ν�tAa ��ը�*�|�IO2�%�ѱ���}0�K�Shl��@?/�����֝e�,F��������{ݍ>:*G��� ����[^4=�P��U���d%z��5��@/TBˠ �����%)L�d��M�lt� =���w�2?�̈&$1VƩRX+,�a��<6E߶{�h�
GG�ӚnN�|�`��`�H�F�(F�����J���o/;9�����a]��7W�#�������JC��W�C��D�����_��%��=f����D�M��>���:F\�r����]� 7�\�v���r���sЫ�;��*�#����y��U�UU���"???�63�lYK˛�c(K�����?|��ԣi扄���=VTU��ؠqw�o��~:�-c��b����6�������!��k+�4�h3�|7�M�C����,����5��l��C���I���J��ɼ�|k�}0�6N%L���i��\����L���P����7���ia���Ðe t�����-�O�(/P�8p�6,�t����[�D)Q}���*��ޤ�3n�>�]]7.E��yg(��ڒ6��uV$�����U:��z��lPx��כ �Q��Հ/���c���O-|�v�4~�݉�a����N�W_��!�ܹ����?v��)�M͂7�Y��1��R�:%�~�S�}˴î-��PK�qW}��B�p��nS:�� �=8���%`yP�{�d�� �vb���X���{Ga���$��d��ՈG2KY����h�Q�ȯ����uQ��؎�0�l�c;L�[>R����=ZM���|�L{�=��յ�����x>���&I���f"�����vgwR��I���曒YV+XVA�Ap�F��SB���G�q�5��z~I���뜺L��À��1G�%000__�3MDOo��-��w{zEEs'>����p,BZ_���3OL{�T3��5%�J��!�����:��E>{y_��`H\G[5�>"Q��h�{��!/�l��w�n��}\�嚱���k8e�Z��Ύ���忥�+�U"���

0��q���zv��(:J#��c?o%"}��[����>�`Et����u=+^�����1_jO��D_O��LF
7~A��}�'��fDDFV��+O;�t͡&�i T�r��LӉ��V�gCv�pՉ3��+�펙u_�^�<��W٭��T�T�J�7qŨ��)_^P�����L����<)׷��M��R�\�������)' ,`�^��&�T�N���B��8�1nK���,ů�Cs!Qp�a�K���Q�6gL 
���VA8��g7}�����Ľ�:�5�bdp��-;*n�ɶ��ib�}o��P�q��|���`����W�*��>2��8�~�E�a�q�+�+�ݣ�_�����7m�w�Y�O����A���I�iy*BuFpxlL��Q{��MV��d䅔�T��Tm8����R&3J-��N���VaD�@WwwEU��2���:{�{��8q˄�~�}� ���G|���^lb%C׬���a=�y��I�++���B$�H������<�g0��R����h���uT�|����FZ��b۷����E�0?V����r�no[$���SH�ˊ�����s6tZ������x�K��>>��='}��

nn7�b�Ġ�����������[
뗉^U���6O�X�cŮP�����Z�_�
�ۜl'��v����7�~�!��:K�I�"�!KsF�7t��..9��=q�G>Պ߿A;]�&u�E�Ҳ�����g�Oy�^���0����zA�t�t�}�����L�?
5��AJZZ�f�%2�� ��j��e�7ݳ��)وL�߆����΄W�=�����8+++�X���`����G+77	d'������)C�?++�����M�,E��~̓�V�.���o`���U��u�^�Q7p���������Q�k浇˾�/e����Xp�	��P *M�M���>��^��[lS�SBO"��	���L��3�O�:aa������:---�	T��~��g�&�9� �'�q�-*Z�y( ��O�o�R-'!%������f��8�c�4����c:>y�A�G�����e�
a"T�!ST��G������A]==s�]S�~p����{{{��" ���2@��;�\`����:vj��ҡ�pq=�ڜ����Bo+?{�c�P���q��9$L.W�Ȝ�g�Y���Wou�������Ւ--��(Ym�e!��,c��F����졲�J�&T���(d�R�&&��3s?��������ݯs���z/׹�G^O���sD���9��E�.�*�O�3\�V��j��Մ���历_�UQ���K���+��V��������ˎ,{���_=��E�/�QTT_YY��Rl�Pﳼ�jv)x?����D1�~�/�W*Y\<���7%����22�~�2����4����'Ѿ
���0�&��9�2�߅���-3M���]z�)�]V{3'�{{꫰��-Y�9��ⶀJ��K�.��R鶰��r�2 T�^��	}���k���� 9>����a�O]ll����A���ꔕy%�����_��[�{���Xp� ,��t�S�2y�-���,��]ua���}�m�����r�b<��B�{��Tx�W�_�q))))��w�}Ꝭ�m`�+W��}9^SS����C�g�����|~{;*+����|����?:%�+vra����T!#&JO��������
H��
�ujW�*]�P��+�Y2�p�.}~^9����73���0�qQ�"��ߔ��|�/E,���'���c���=����A7;�+m�I����"��::��{S��K���k:�(^��+���U��4|��S�@���:�;^7�����p��>qږim�{Ğs�Xj�aƥ����ɫ��I����Kbmdd�Y��`��������hЮ<�oh�������5O������?bt]�,LP����q��k�+�]�2	��rͣ= u�!���ӝ��,i�M������
�v��y�i��޸Z��ձ5�HH��-.$�z�3o	*�E X���.�������Ӄ�怷�#T(�**Y��K��꒢�֙��vZ��� QN�������}��?�޶�6���ގ�Ћw���KAA��ӳ�/��MLL��[���q��2��銊�#C�N���nh��\"��{�fq��1i��;-������͵SE�Q������O�������_^W�"'��[ZjUj�p�MѨ����f��yiiihK�b=$Q��H��
�DM3s�?�72!c���'��2ԗ��@|���OmҸ�066l�5%���f�Bw���e+���5qў|g&= µ5�?XKѡP(��5�o�!�����ymx�p��l$�Ç�FG�8��GG/�$ܸ���V�d�z��ŧ ��b��*�"�Κ;��;Y$r�n�s��#�����z��ŋw��U׉%�u�%z�&|���;32�]3��6�[d��CX#��D$H�۷o���.�+�,����;Z��(P�wv��Z�5���ɯ_� jÂ_�|��5�p�۷m�&Qs�*��<73CJ�=��4�ɨ�S}�߭}!))�� �o�Q�}��1�Sh�o�^�ݽ������Ҿ``o'?�3�a	��?��e��l-v0]���|�Ȧ��@x
N(�!��v�`X������
>![�}=:%���nm}xK��L&������L�=�������	���Nb8����Ƈ���3�Vig��qx������,0�

�CC�0Ň���A����E?C�.�з��|�&s&�����D�=B1��4{��s�LDf9X?:�<�/��h��t��@j�0�,�iei_��終ώ�<���Ó'������M�|��u��09�ap��	Ԣ<��87�����G�\R�UQ]]ޔ�'��hk;�Yk=V��NGG��ԛ�R8�����@�������� �[s�G!�Ү�@F�FrF���!��x��7T���ҩ_� �=L��!z����V��I�^Z2xQPV�>�U8.s�n�ؾ��0�ea��O��+�k��]�|ܺ�r��M�ߥ��Ӱ���w��"�t۸O���M��C�2��
�k���(ͨ:������V��`p�"�_Ł�{�Aw]��vq��}.q��e/�`��,oHw�X�M �f���1v}HU�zWV2�lٲc���	��))�9D�bEE�#5�K}��Ve��Ь_@J���ˬ}n�"-b��vf)R��)5F�W�Ė𻜪�T�t����__Z^���Br�Qi��c�kA�����h��

K>k�R���atj!#�4q��!9ע��J�By,�|�=��x�&
����Ԕ�W��J���J���[��S^GmB���h�]����Ꙓ��{���©���:��~������������쑻��`R�{Ǩ���@��S�ڟ���li���R::n��t`�c�� �Tq����]���&k�Vʘô��ZYY1nsb�h�/�#��`>'k��+"ӿ���o�){[Ў�!<TH�s�����)W\W���n,�ݘW�=�V=H@��S2,��	� �<�L1���AKED�uu�u�����q2)D[V��O/L��t6����EG�J�j����{D�^��KJv�)w�L�0�4j3O޵�*��Y(S�{��;:���ז������6�6�B`��jk�z�vlD}*���#�-
Y�f�=C?@����uk� �\+�L��C4;�U�6`_���65|���!�w
��Q1w8��{(D�b�L�T���[�0LQv�� |�!e��5c6��t�4�5���yy=Q��Hyd�<�߭T^����7���5s��^p��|��D��kW<�:���p��UL��O��~����穽;7�C�D"m�\��J�E����d�ě��~z��L�4�ş�����ǌ�|�߈�SZ��yә ��Tb����@S��]�9�W�Rk��WU/0��4鉠pɕ�G�w�|�j��/��:(0���̚�qg�g��g�m7�a��X�%�5ƵĞ�ޔ�?i��&󨝡Lˏ�y�v�)�@r������5Sy*������<<�?���}�f�/��Z�����ξ.��;�@�?T���n������y
f�/�eW������g�m��K�C�>.++C���С����������ʸ��6%���d�t����P���jo=$�h���=F��X%_��1Q=~&����a�������k�d�`.6U�^d���ݎ�svt<������TESS��ݷX���+`bll���+e<K��ikw@J��\��G�@vddCj�+�Ϡ�g�Ev1�t^�"��j�ݨ.�Շׯ�AG��=MJ�(GT'�����>���s	�		����$n���`�+�3X^^���7\H8^�����,wQ��@�#:W����ݭ�<�;��\^�����ޓYz���J[�K].��B�Đ��/J5�L6i�.7O_����K8���Ŀ>;/"�J-a�A�}�Bz�ϴ����Ctt��W�u����=�A bl��ӂ!�]��@>�U���!A����)������1�}6{LZ:�'�i�a˵Hc/���B@x���g��<�e�W�d�V�}�n����_�E��ߌ�p���FAnL��!?�=1���$:.�#��^�{К[,�}bb�Drr2D<�$�fvv���t��HN��ڝ�||�R2ݻg�� |;6�t��7�fm�XF�쬀�nW������� X�o��c2j^qB=�sq��<Wa����������r��q[*jj�XXtoڙ�^�	G��%�%v�"�������>H�������+���5��MMi�~ yq8��dgg����±b�.jycc!�H|�.�D��{�d]˗P�@
**�4y��s��^f�F����J�v�i�s�U��Ó7Ng.8�SVV�+F`ejzA��%e�0��b�d���-,-�&&�d��/���H���� |,l
{�C����	��wM��?���tO���6E�]��	c����O����V����O$��~k(-z�[÷�e�	�y;��o7uD�[�=b��fV�<�'P�B�Y�Q8��������������ń��/ttt|����.&{��,.���xT�~(�}G��}!�*G�Z;���)*�d7>a��oĕ��E���̻*?��P%G2[� �-ZP1��}t��E�I�A�D�-�Ʌ���#������d�=�aO\�aXX��̔O�^��ȫ���^	����;�NM�*�`�r�n�gd譴&$����)"MAV9Y~�� ��_��"-�����\�<�ڂ�a)hz��)�LFG���SDFN��sDD�ĸ�qEg�V�թ�隁 >}����w��<o<�������z�������6sPt\���$��X�剠=��L��_�jt�>Ä�K�;s�L���d�,lXEʃ���E6��uu����M�#�[�����L }J#^���8�rkhA�ð�N� �z?[�q���

f����5��o�?�:�se�kj�b)O)�I'����$�jӹ����J�[���D-��>)��7�#����t��&?F�ۭ��r�9����W;���q�������,r� �9����skFx��I���/��5,M�
���LO����ֿ�Y������� 9Y٧���)���T [*՛_@@4�!�p��T:rĜڥ�诗�)!?r���VVBo��F uAt v~f���E|�^MZ��3>o2��8	wx�P�腀�]؇^t��$���l��5��8�dť��@||��ܻ�x��w�2����h�����ݳ��J���[�5�z''ol��0K��|t���jˆ���ٌ�ޚ���#;���1�SS��q��ZG�3�**v����nn����̨D:�Y?�ևd����0��\-D��]�#�f��\K����XU%rcC��$.G_Qe��	�_����m}��5^n��E�xo6���G�Ch���z���Գ�M���::;�_<M����7JԬAz�ZAa[jZZ)�D�ڜ;������heȆ�mш�+��C�.��m���fF� �k��'������ͨ��sX�7�5�y���߾��vC���O,�0ͼ��:L��\�q?7�!�H��������6��:��5��J$t��W�ъA���F�r���o�v9�����J$&0n_IU��ř�!�'���LH[�D�XI�|ӦR�Tb�{yUU����jH�e4���*�tJ��qb|�
��WS.n�=59�T���9C+$��� |��a?�`
0 �D$�[u�-�2���P��Ӎ�Oʹ2ܷ�	�korj٥	8�~�bOb�^�����N��j��G��J>�%�����ڇ�w�UgeYC��ޝx:]C{����nU�n,<Y4��'x��llc���,,�@�>!MHެ�����r� ���͑�ԓ����岪�� �@�����n���Z�;I�]td��1��ە��8��i�����埓�Ew���3WH�_?F��)z
�~��������G��
��/xB�u�n̿�w޿m!�W�����)馼/@/���ܕꔚ��A7�+\ve�Z��C$yAډ�cJq;l$��3%*=G73�;��"� �	�jɐ��)�����#��tB�����l��]s?kj�	d� �A�W�N��,`��D�@�E����Vk��p�"���I�7T�WL��?U[��t�����=����'�v=��u�|��>`�9�H+{�z��^G����Js�4Nt�څcF�>�z�x@�3@����h���!y��v�����o ^Ss���QAQq:t�y�y���
��:~nYi.|`&d�E��BC1���J7{{cF7u�8��b�yA$\��G����,�6���Y^F@���<r:���(s	�����5)��,҇������Nn�k����2���V`H!e`�w�И
}7a��1�f�Sp##6VV=�O� ����|��,++nh���c@fQr��T��׮�G��i+�?��{V����i�t]���Jim��ٹ������7�9!~�RߠB6�ÚC��sO>޸��Ѧ���������z�({㶤{k�Xo:�6��7$��ܢ2�A����{O��$��-a9X�BJ��h;R:GwA�0������P3I3�x��rN�;��gf�7]g:A��`r���]J���_2\co�599�d$V�����Oo=_6��p�v�����/I�\޾��ƙo�jPaֳ��M��>pxG���d�\��1;��Х��ߜ�XN��\�066�;l\;XRY�bĹ֪�S���=wA*����W��oE�*3�}����r��4�$50#�o�Ĥ�z�/9 �c^�`Z�	ߙ�zQW�<�����RJII�0E�&���H����V�-z�O��L݀4ٱ6tt�j\����۠rf`�Zh~avP����K�pkg1�D<���~��ZQT���%���gYJ#�ޱ%Ŏ�o�j+rC�.n}��ME6lx���{�S�AV	�]-'�uSN��Oт�F��ԏ�)%d{�6t�a�	v���L%����'��)��C���r㢽�������s�4���KP��2�y��qE8���DF�Ȭ��^���w��?�V@r<P��`�*~c(��N���]�P�Ha���Z��ZG�i���u��l_[	�eb�0�D��c|ㅖ�E����Ś�L�
,�ȹ�Y Ƛ�"����p���q�s�"�g��!��cW���P��d-kC ҿgOk�D���������~~��IZ�Yu,`�v[�,1F������2�6�u�̟Ǖܻ��:��B\�Br��I�G��ϮW:�2�󖽽D8,,�Z�F!���׸n��+�i쁥�-�(Q��� }ĭ�4] �[���z�V�%w�Rː�Z��l\*����kᓱ��g����96�|�%����ŏ6X<�E���l�/�]-+sY��Z>oh�*O[φ���kR������ʪ����=�X32.���+�M��*ͫ�2+ޓΆI�ɤ����L�� Za��W�����f�10�P^�P���s�E�U����ʔ�e~!���a�Ɯ�!���k��9g���̔��5Ct�(��Ҹ ���[Nf��=_��Í�6]Q�"���#UC�huMv%e��(�Q��-���Y�w>*�B����Srs�C͢N^�:�?VfY�g6cX�����=7w����Ϳ��F�
�K���ۂE��rso�������77�k��L��1����L)��]�h��7�C��o�ml�7����O��p���9�fiQb����v�.ګ�`"�h7�}�&�&z����75S��<:�a����>�7[�����|�5Kˍ���Z�m�S>�.2� 5t7ĻU�������\f��K:v�chu\P@�}MC@>���׶��dz�����0�+����+gV	��0�W�mҸC��Nx��]�^�����.��^&�u�Ndۍ��b�8�@t/;*"� B@����i��g�b�=u�w2P�N�Wl�tK�\YQ[���DY'�S�rqp8c�v0 SR��v���&��gx���Rj;=6M��6�`��1#�0�q&j�F�rei4�Ce�C���(����Ak*�̦�Q�_�}��Z��C���6+���bî��%?�h���>+L�ܔO!i��Aw�s T�8��X)���_Dݚ��n��N���3S�!���:�hr�mr^���O2��͘6�,��~�X�y;Gkk5���3V�.Mt����z`�>f`�s���X7)}�^�	�4 =����P��)9T��gJ��U���֞�!�S��t	UCh�e�n*����E&���u���3ƝƋ����E}�a�j
ƶFi�߭�������V�f�Я;7`φ^I������wz�T�o���?�5_<�o��E/G&hΦE���G0�C��ֹ��e`^y�2K��":��q5�����\��:5�n�5�@��1/�wc�rr��_��q6���]+==R���{�ď[n��NMJJN����h�^=��<��2Ǳ������C{��q�}2�m�r-���ʦ���T٫�cHe�m�+w�k�0��#0���7n�)J���3�*���;8�F-"Ħs���r/o����hȭ��.����~N[w<���>a�6��)io��I2*%�C-�#4��w����l��j�@ ���-&{j{޳�[�qnra��bߘ|真��C�J�1�ƛOi!��7���F]\\D�q�W�)us�ҞI��;[��p-z��0�C}�D����IY@�����M疖�����8�2S���r��i��=��8�D }�T�פ U������;ZVV��\��se�:�A`����<�>�M�V$�-������"_*���}B�@Ƭ@�!�vG�$j:ySo�~j��q���ő��+�l��.��HOTe���+ �c�����aG���u�a%��u}����믕�S��B�DE7��I�'��.]
�pJ��A��r��$v��W�SqII�t~����/3@�[8�S |��0\�M��*|�n�J�cY���.�`�ii� �_^~�Xp�ā�5V]�ڰj����uto}�|y��[TjG��TZmm�>��U	,��ELh"aLV.�@29aD~�bX�`�b �]�6��e�:��P��y��ϕ0�@�ܜ��񮾚�ӻ�m�ҧ��{񌾝g76 �p�ڥ.s���;�ZfV�a����lR^^�����b��d�9C0��kj.��RK�K=��i�ZQ�����WKU�.��E��/$��LT��/��~"+�B��Z@/�8��[�JKKKM}K��㓟�^5���9�^�m���O����v���U��S폱G��ۻ��sF]S���4�4ݹ�.�Q(F2Zt��Op�%)�Xi��kf[й�v�E	�@�Rף�����ܫ�Y�C�=�u�N�1�
�K�4�AG.4-'�!�zN�88��?�dK�~Jȇ\\�Q�o��`���3>|�&n�����s"CxLsi�Do���`��E'ｉ�}�d;���|����	���J;�'�!*QG�l��������Հ���Fy�S;�uܧm� Ϙ�u�4��= R&��{�%�WF����&)ɫ������e韸��S�v��U���ң��. ��<��3p�x��5] �\�|�6��D�iiy�؅�mQ��wv��u�$��qT�K��A�q�%���?��y���08G�(SwZ믤����!@|���b1T�;?P3N��K��9��1��S܊C�xMmu�����
��q,J�5J��6��Ӛ��q��;q7�hGSN�r��&\��'���4��^&1ݵظ�v�y67#��r&�{�P�m����ڔ7u�u����l1Ցv�����C�.������1~�/�:$�*<�FY��d��k����g�v���>|���,V��<G���7�5& i�j��8�-�}��ݘ�Bc_����iŝ,������ݗT�}�0$����^<�Z�x �8Chp�0(Ez�9�,�h+�ZLzH,�fo���Z���;WVyP�����v`��#���R ��VK6]���w�0��u.�q���� 	oC`�{�f�$!������<���twOO"D��l'Q���c,��!��`[a�9�.���:�1ݘy�dB����&$���RrM7G\>�-��]�g���}��f�����x^�S�X�*���=lڷ�������d���ʚ�/$`BL� ��>��J��,1+>_av��l��זa�'S�?9 "�q�\�`�fk�A�z�Y��,/
�1��q��;�����UU/�	
���h<��4����6W�A�'|��]�D��`�7R�b��&h����x�L[n���g���j���]}�"�����*@7�����>���4��:�Jd7��n������
ћkl�젛z�Tk���i!۶�����K���;�x�U
��M�$����7.%��(J�C\�i�Fu�����c��%���܍nd�d��-���d�[�G�Ú�HOc�Ʉ1�R�>��jm�ҴB�	���Xp"�ԧ�Wt��r��Ҧ�A�����E=�E����9�d��������r|���$/���ri\0iH��{;��o������C4��<�Ǹ(gf�\����2��w��V�Q��
khr�6n� @J���k`���r'AX�@��I�9?�O�YZz)R|�w���Gx)Xt�'������(�$��E^�%"���[�U��9��[t+��F33c�:U�[潉}���ht϶5o�M�clB��4��_Z���}����kB�oO���O�-|�p�����y��l�{���}��@�6_�5rP�w"�5���99cl:֛���~Ϙo^�.o�T|�}J}R9-����g�R��G�:yԨ3M�XE^���s*��ey���l��s�M�=P�2(�/f�8H��ĭ�%��	0^� ����:���;��ew��˩����&��5�8h\��6#W������VC����La%�kgJn�+}hb��D���C332�<�'�~i�)��c�*e��(��=��X�^p�m��q�۱���5�� H+���>
W��V�O�������N&��}m�0|������4d��n`C�1����Ae.���q�2s:=�$ȭ�o�B�3�!r��3�w�A�,-R��Mpe��=�o�9���3ss���'�85ni�a
l�2��K�d��h�({[t����Ύ���E�@���^W�1�5������
�Y�by��rG;W��+$= �ܢ�XƩ��y�YX�x��죀zL&��U��͗_p����?�щ󀇰��q�\��<���������sv_h�t��>���,lP�q�D�S��8$���+���N��>x�;��A�AW{�]s��e����T���d��J�ߡ9��:�q�
�v|�����ƻ�A��S����6��Yw�:�ͦ���^  ڊ
|q�����׏291q�Ҏ����637'uJΊ�L}����F��ٿG�CW;� ��
�gE��P�V(���Wң���v@���	fffIN��كt!PV&���y{�-����2��`�
�3!��4z���!t%�r쟋IŶ2�5m�k˵�3�d~Y����yW�h������ҟ�h��F�sC3o�V��d4��5=�\�%Zsgٙ6���<O7|^��$�\�\F�(�d������d��Ø��O���~�T���}�f����Fx�};�����nP�D�@�M!v��s���/�kγ.��q�;��E�!��4��4�.�(���w9��'�Pҝ����#�s��<�:PL\�H,�A��L�o!��)ߺ�X��1����'g$�6�����M�g�%�wSb�'�~�V��o��
�u8�����lsj}�����G&�=��<A��-7G��`�ڗg(l^��.� .yqCa+}�y��q{�ν��ۿ-3$t�������A݌ǀ �V�;�K�ݭ~P�#��b~����w��_��,/��qQ�b�M2������<Ig^�Zp�`��lN2KZ�n�[�¤wf][��9��ZO��x�B=Qx�����q'��΀�hH���	P�Y����(�����Z-K������������;�*w%��TZ��m�u]�P��-�R��4�����i�����չc�k�ux~|]z�p�9p��۰����II���~y�����x#�5�e�v��qp#' �ε�*��`=<,\ȿu�2h�L'^���<um�^⋧� z���;b(�\��Xb(���?������S~�oqG�kٟ���:�+�˕�h�4��t�!�gȜ:�JYWCײ7�c��!t����D�8��uj���N�� �v���n�7�H�*;�U�0�� )ɮu�t�8	�_eG�bz%���S����㲣�N��|�B�b5e�ŏ�0���r�; jb����n��ә��Fe��
DY+6�ymϜ��	9���f�q`sD�I�u��AjzzO*�ȏG�`?~�����h���,J\P�Q4ں?�b;��&k	 kq��e�Ly,�Er���_	\��2)s�o2�����������_K�#�9�#�K���p���S���j$�<�y�:|�*���9KP��� �h���vU��׮ᓚkC�Q�?���J t������1�W.r]�^i�!B��oD$�ġC�\��Ls�T�n��U�e���� ��fN��E�V^�j�D��~�5V���&�����oZM4c����+A��>��)*Y����Ό&��0�X�V# A��|w�3�%@��Ж37��Iڂ�3o�֞�����y��Y�k�-�ί�P}rle�3O5|	����u���9끭,J� 8}}u���9G��(4.��!Ϥe�(7����?���J��Z��芠����:{����0�A`7�؉��B�Vu���H�Ufe��հ\��24s�;�xv�j�������o�)M�� \��]e.D�Y���,�Nf�iiğ?on����s:;��Ԕ�+�ڿ��x��������]��S�//�s���rϟ]�$��ӕ�����rU���	�4�ي�G��--��X��be����z�w�����o�fΧc�J��@�x /�$v:R�
�-l^��Ҡ{�b"v�!3�����o�����mm=��$6lW-YU*�Lh��ts�� �5`(�8㤩9��Z���@�}��� 
�Ʒ�A��!���wa�-�4�WwG�����]��g�7�Vڟgi�����!������!3C�!�ˡM]sb�^;�o17f�m���(�5Ue��V����V�n.�v@޼>�!}U�J�[Tw����G�Ywh�����4GF$yB�V����C9�aa� ���X�ΑN�^k���F��+�L+]��-���<���T��F�.�h ��|��>ey��1�ԑ#;���5U�3-K��cϵHߒރ��A���Y�'���++-�H�C���3M�C��ۏ̪�qO�����
a����m�7^݁Ef"SYE�y�B�O��i��ο/�X��5�?��c�wÚ�-58�Z�B��E�t��`Q�
�vʗ���N��fo�\{����ǆb�! $���D1��,�.r@a��A��d�|�zUI�[�Z����^����1���[�{�K�5�������]���A0=����f�W��J�3�I��ip�-�]�.���d�RZ�R��j���FQ��k���u��ČP��T%K����z��\�DS�h�-�ٛk1??w��Ѵۊ�>��AyT*���M����S�����<5N��e6�y�w��ø��'OF�+�^��b?
�K�I9}}�I���=��/H�w���a�Af�"A���JlWzcB�1�D5�|�0m���(c�gc��
�]��.̟�����Sc�ĳJ���F�)tE��5����|m_�z�k�.Ձ�#{.�zVVZ}����2)Z�M:��؆�'��|)/��[sdRY���9H�U�h��uX��\�B�(�s֫=r^�@�Hs���0����_��α5퍤->��/4��){���s��c���x��C��Z�#4����Z��'��)�*��sd4�]� M �ǋ��X?"��'5p��.�������.�[$퇒ILw��X��U���Z�\�\W���0^�J�_<"�D�fr3ƾ,�̢�����]����� �{ᅬjӣ������������11)~�)���v[d�S@��|�pXj,������V�6��Ufwth��C�N���N�����U98(#���a���6^6t%��c�&
��$wvv�&/�i��>8��ЛkJ��&{�f  ���n������Ǭ�h�����ކF��Y	�Rf0e5�^���J=�����Hk�ng\r������my�M�'����B_"���B���J�⇗/Q�i�p�Z,�FC����Ds� M�U�C��0��$�������VW?��R7��W����Ӄ����M;c� �%��i�5�m��ݞ������p������a����Ԇ�����@�y#~<n;��񀌡��b�R?���M��I��8ŸS�l�J�cP�]ӓ��(k����[ɹ���^�@}�~��L�<2��.�%v[��ac�+���s�ݺm��D]G�J7��ס��C�bMJ��^�2�	��������5�e�����d\�y���(=?$"�g�9Y9��TD����}<_���W��r�J3I�j�ݭ��A�'''W��i��{�T�UMi��*G�`��n�����4�Y������ik�	��._

���u@�������m��\~NMi�����d��<q��tq�f��A�jN��n�uJ�z����� ��O�����7N
Ƞ�Zs�x�~;WsI��yq�����>�)��r���������v%	�ր*	\����M���֞�Y�Q==��"}	��r�'3���J�nd�4}�jC��q��0<�f"�D�A���m\��rǿD��� 99vv2)g�H�rg�$�Ҷ>ał�`q��z�P�Y?�+(tO:-�⣭�&مď�y3I��d#�D�c-�^)������l+Ã��}�ωce��vn����]�o�����t�����n]T!��Ҹh�9��kg�~��6~V M~���N�[<���c�0�����h��e�����(u3�(��������������([�ͨfT���Ie�[������R�m���l����!��n �ԅZ��*�F��!��\ߢ�������g�a.E@CӤ�>S��xJ��Q��nk�5�"��]z*��QQ�wƶ���V����?ɸ�q�6��u��[�P��8} Q<��Hգyx�;������j7F�Fe�#G� H�
�v�~"���J���Ξ��
�>�����f\5N�;�0�Q��V��W�{�A���Y�BY}�\��ˢ�����g�y�W�ä$c�NP��Dp���[�0�̏��ԋ%��"�
�7`��ϲa՛Z�Qsr2
9��p��P�A���;(�9�h7��[���~�n�Z�1�]���^av�_P���X��/�6T��.4srw�\�;B�3'�3@���y`��- U{z���ڭ�뎁PI�y�)����\P��c��3��RJ��J�g�^$!�D�ؓ�iugD>~���dT$*Ǥ�+�5���=���b<�qnrtTz�Fߺo-6cg�����10A�R�U\"5 �k
>�/���p�����$�M��\{�p�am����P!���/�xoo�}̷T���
�5`$�L����7��C�w�2D�ls��)��Vq#�!!�>
���_jY�{/K�ڙ*6΅	߰z���<�j��61x�Z�㌧֍�ي�Sb��޾��V��d�TԄ���֩M�b�������\��h�.|uǺ�L�κ}u&{�y�����[Ǵ�`C'��PG��c2���2Vӟ��$�ס��}�P��lǙ�q�u�E�c�zn2V����ܱc���IvʁMB�E=>>>�
���:.��q#�a�gM�=֪=�����o�B&t0]Gj��^��0��*�U������/0������!�lSB0D���$�!�
�	��CV/K�U>��r��ZL�st�Io�Q���C��ds@DE���N4���|D�1�5��߆��`���
5۴�<�����k�M-A��Q��A��a��:%E�֮;� Fǹ#�z_<�TrZ�w����e#�>�����l�㲓���7Q(j�zg;����(��7��C�X�	���1�����Nv#�n���7�rF���^��"مn��h��B!�r)�\?���������\�Ʒ[�^C���m]7L�,�Gd������� x����8v�C�9\�k�����	����ǐ�Z����9�碷v��q�l�֣u� �y��Um3�)��b 0��-U�U�4�G���p��ZV�@$�H��� f��Oy�|[�X؃�.=��}�m:������.0{l�.�˥������c���d�36�:�1�-]R���b�Je�`�z܌�`k6��7N�)��^�э�������Oh��� i�:c�Z5: �k�4N[�)�W`0*"c��L��˗*\�4ow`�k�)+�����s���}zB��I����	w�y��|^N��7R��o��,k� ��U�tqq�a2	�Vh\�p������}������m�D|}����R��.^�0��n.nn���v��u��i?S^�8�G<����w�R'�_`:s��a~~����?`eE�<��UD�"�" ��OP|�����69vv͉.�aQ:�蛘\���F�ȃ�2K�S�����%jLd������C�0���s�r&�@f[:+`�w�f�=��;7��9m(��|Tʨ8c�W�x�~.�4�s�[� 7�~���>���?|Bt*.�8�U��' ���/7�
�㕠��7J̋�ኚ��A80̥�	�:�②,��4�[Xs��<3�~7���>W��B� ͝;�t��88-����+�p\�e#�g�B��Aki�F��㘃=s�7�QbQ	i������Dͱ�y�[ֳ�8�At���KF�K�Ҳ�=r$[���M���~��k<�F��1*q�2��c�n��ݳ uԙ�[��w�:�`g�I[Gg�'��%X�(�O��W�i���M-ޝ� �Xt�W��K�����WP]܄�c@x �#qפ<�����]W�p�Q���cF!@���5�.| @"Q�T.ϘY].-��X�'�,q���1�5�T�]�anF�;��_�f��Q�Qz&)�w&n����&��kzl��[�8��w෕3M������3���06�ç��f�K�b�B�B���P|�N���Rƅ��۝
`��v������ �=�	��:��j|c��߃.,^e�OP|����Y�&��M�S�!�.��H�B� ��>sB�ݎ�(m�?}c�%D�M��B/?K�5�}B�(2+΅�;�|j`�~x�qqٝ���u��!�f@��e�/���þp�;@�g0�-���4��/�[\�#4��x)�XѨ�؀�~�|�q)bz���ʹJ~����Sx�u�-ҟ�Y0]u��KK��\{y!Hbb茰����Ў̡�!�I��n(���#���B����'��`�:J�ŚW��}�0���9���#Gv�%��s�?A	/<$������qvsS��&�r��o�f`�T=�L�?s��0�1x�b��~�Z`%�������hJ�K)��v��5]����u?��(@��.?�,ݽ���!P,�Δ\Ђ�7��@'2��SÇz
����	T�� �~�����[�\��k��'���X,�?Q�"Y�L8�7 �p���Vp�LD3��f��>9<�9�;��4W��#�L)�Qƕ��1�j��-�k���4s��#���L�2�����֌"*c#
�q#�$X�Qy��q�0;
��55�M\�,��q�����M��L�������;{5�D1����ʨ�	���H$�!�TNO��X�2�����oYZ`YJ��E�k���qS,Q�x�tB��=...�bX�vZ�)�%	Bo-hƑ��ҫ]^t�gU��k��\�/���A���HT��\��\qu�Z���a>�J��I�.p牡X�ҕ�ݔ��o9�RYyq�ѷ�k�H@�_&A�+H�$�eV
-,r�;�"�i0Op����� .�����s,K� :�f;�E�<��II�PNٕ��I��WĆc!@kڒ}.��=^�8��y<�x��Q]�\�E��dŏ>[�/n$_�;���b���K�z��z���Gd=d�_3�&�
�eR�>�@������`�ް'��?���B�Ƭ�2�X�����ፆ>ˌ�����յj��u��kԧ�

�¨4��q��	��^���p$�r��<���~�J�!���r��IT�ރ���OF;�ŸЌ�b�*������Nˤ��d.I+��c���U/��f�3�2s	�ڨ�Ь���"�8ϛ����{��@~M�֩+r`� 3BQjFR�Ad+�0����2��`�?R�=�-���V� "X,777:����GT�7�x���h�,�p�ϕ|�quA/K�P�.�Ԣ���QQ:�_���K�&]�|��n�W����=X���$�1�ƘC��Ы�F�p�y�� �.��E��9fm����B����yfI�b�U0,Z$�=_OT,S�10�,�p} �_=gUE48�Mx�~�Pnn6\V_<ѫ3����P�v�p���G�C��!!F��S8�@/�CȰ��-�NT��zL���1�`fON���$������XA��_8d������u	���y��f�9�]#S��v���_e�!ͼ���0��N�8u y��w�j��CѸ��r>�D|�E%&�}zFy&]A��Ȳt���K�ܸ�`x��K_��2p�jlKKH�s7��ǻ���^9[���cm(└�aP:��C��E�.��Z[�����������j�����&�P�o��t:'�ꤨ,�RT
5!kG!Ր4��![�]�%ˉP�J��,�ݠ��11֡���`01��~����_�N�>��<�}_�u]�������ۗ�((8�δw,4=�.��=��$�\|y{g�e����a�O���0c{�%�x�,F�Ըs$��E���R�l��W�Q����r��������O-��|�����zi��\�ḟϟZ�{A�˵J�.���ik������s���@E�n@gS�t�`t�@!X� ����Ǜ�C�y��⪗[�)�feC�-S�j܏홥.}=5�D�rd�:�͛����_7�;R�)���%u��Ⱦ�~����pW����R�"�<sl�`{:�M�����WV<O7 r+�vt;�̨p�|r{AW���V~��SSץe���־P=>,���ޞ�5<-���-OR](�f6-���۷����	�R_�1{�X��7��_nJ5^�>�Ӯ���J��<�3�+������<#�evzl7��@W�69�G���70p:F������e����Z��h�����1����rr�룭ee'�O���SPg�ٯ��

f����������w��XwQWA����|�FK�6�%=���B�F9�Q���{�[�,#�Y]�o@ա ��=~���D�/>���V�����]R"�����$�v�;,~�|�Xh��3t���6��i�'A�fG�g�K������sↂ٪<I�%QI��Q���V<�����Cm�4�\t�� �[��i���R�tH MW�WB���5�C�j��.|ln֌m�.r���8jh$^����ء���ľ}�RS>����S�G�e�L&�������)
�*X�'��w��f��)Hצ���j�������4N�c9�[��xI�!4���b��,L;��u�ķ+�/�?z�YN�۳����pp���VffG�u�Msc[�t1GG��%e=�����a�U�p�&�m�̭Z��õȘP)�:���9))	��?�,[����(�R-���fJ7.q�r��9ʸ��vv����m���1�����^[���Zt}�����pެ
eؚl+(�SW_�~8[�O~�������v�e������Z�~[qu��އ����K3�ns��?�u��b(���Ņ1���hsf雛��,f�v0����g!�j�"�k���###���ή�.��t����IMYy�C�_}s�����a:���	K������ݾ��a�_�md�#ި��Yd�Ht���8��_9���Y�y4m�T�~�&��J��x����(����w�;$�������=���[B�ޟ6����騘��`��zT}��61.�W�CrHV8q.׽��ͷ�\���=�`�-i��9X�dޢ2�A�|!��(A�R���Ɓ��Wx5p���npf�N�pi�:1��?�z��4�[;<�YO���E��Ix��xD`���S�p��kGr��|�2|�x�Kk��77��n�*���5����NjN��P�/�	�<�4&������u_�^��.6��w�[YXD���wvG75e߽���K��^S`ЕV��a_�����z�����l���@ʰ���6-]*<�@�-�y����� �>�6��|�H�R��iK˘��8��	(�2���٬�q5�[�'--���"s*��|���e�Q���[;?_�����G�~�C����P�Z��yʱOK?'c�Ύ�e��4�طhƔ��o���R��Pz�c�$��Q�W�� bup�a���2�C�5Y�)r.���崲��
boedd<c�=�5���7�v�Z�А:&,�Mv,���~HRrr����Ǐ���-NmF���h�[�Q�=���r����Cb`���!�)���4��@�q������RY�
�M�n�%8h�n|�eB��sϘ\�����p�.�f|2�tjV������m/Y)�>��g_������cr���K��_O^{�89��oK3�M��܌��6�t{����T�E�����X��|in8�l-�"k������D�zW�3���
7�#!w�،gg�ڶm۬���{u%kQ���R��y�����Z	�?�lYDӂZ��Eg��H�����^����|]6�hhd��=��T��\_U��Ko�Z[�����w��e֣tg�,��|ƹ4�|�e۞"�����ߠ�V�雖�qȉM� �0�:�N$PW8 ��h�L,��ޕ�{�Ïa��:0�f�!R���Ac���Xܥ�
ڭqNDЇE�gV��F�@�ViQ�W	���0���t5.tuN?�JN��@�XC��Y���^׎��2,]������V3�����d��'IrǏo70�� ���[M�R8�����l��ƺ<L�-�WU��P��)��			��+6s��D�IL�%����;�E�=(&��N���>���dCqS/s�����J�?c��sP����֣T:;������������hY���Ϫ����0���Z1ˢ"##o@�y�єS�{rt˖-��L�SU�]^��8���XUmWvJ$q�Hsw��w����2,�Ѕ3�_�t�a�yF�7��7pc�r}���l�zuXfff�
D{zzt���_8�X\�rNw����Q�|=S�z�� �d�d)>R���5���֜V�����k�S���ựE�J�<��*O`��cTaٳ�P�x%�V<�9?�s�+�[B��P��c�j��$�ÞL�8����2:5�B�l��V��k��Uה:KO��?dv�����`�[	^���E��;37�M|���g��[��p/Ǡ�6�������+պ_��2�s�#��e�G@�rG��a�.�AQz�;�A�,c�˩��=J�o[���=Z�һ�t�@�inn��X�RQ^��0s�<�Pl.-���
�D��ϗ��G^^�ܒ�B�
��7|�S.Ek����ˢ����������I&�)�^��aw�SL�Qi	)��C�Wܥ������j.�	��#��
��a�{��ֲ�5n�w���=5���^ӟr�'ME�\�"8}AJ�Q��=E�gr.Ͼ���7�{Esz�L�˾�	�~�1��|���|�C�A�N���ȗ���zs7O\7fT��MO_f�A��sK�烊�V�����Oɖ<Z>H)��TMQ�H�25L���p�L�� ������ĪP�+~s�`ƫ+�g^vwuE�R�lk��R*�� ��B��w*A�����$�5���.�>��� �v��s���e9i)K�`�ҍR�08k�2�������-�3����TmV)+�B/0�, �Ɖ� ����rn��l�0�Eƪ�I&��!���/��N}?�O�9�L���V�4���)a�2*T��*�Lf�����C>��kв���]̡Ξ�)�㣇ɉħ�q�'M�iqd��xƩ��L�j�Rǧy�������.?��fm�*�F�W��p�,�~Y��,#�J]_�\nt4��֒rPjh]�2��΢l&���1xi�f%�(h��w�GHY�T�>�x����2x�\ӂ�2f����n�5���ӟ�j�/.yr���T"IoY%��T��\lU���k�rD�a�N瞺Ky[����Њ����2G�S��p��[@V���cJ�-�B�-{K܃����"�A��}�`��՗`�"������9��p����|�����ԪR߾��O��b~wѽ2�g�ީϕ�+�y��uW�*rN���jf���ܣf��@7�|h�2�:�m��Յ�*��Xڂ�k���,��#�RO�H<��*�k���9_:F�O�3��)�s*����=kI���*(آ���أx�����W	A�QI>�����L��osCc�즞=ل���3�VG�7��I#�=��;�TD�2���!ђv�����XC����/�L�s �a����\���(����s�jn�w������@b��`]$sr���I�#���6�/<�COZ��X��z�������e��B[�;�@�2G�=K�2�[��K�SaÚ� �~J%���a�c�lq���C���ma) w��5���<��p(3�e����=v@k�"�Ƈ����82$Z�h��	m��e���-[Z�1��L]�H$Yؿ[�(����˟kn2����j\�A�����c���LA�F��m/���'��Ř]����D��s�'m4���z7X3���a���[AnچZNY󷵎�C���y��Է3_
������-b^�=YM����y�:{�!_��b���ӜRN�mW\Y������f`8G���2g�e���=	0����9%�)�O��LHS�T.����fw�ݐ����m����q��-� �GOY�,�ฟ��HV_6�b��N撓���e�Db���@�<v?�����{��i @>"1H�XD���qֱ�̭������C�f���e�\)0�K2���_�4$�I�W�xE��ѹ�)�֛B�ۘ �M�����nT3�͸�����2�K��?����-G4��b�`�SNqUK*w)�v�dh�ق�T���6��C�u����*`#X�DhEn��E5��O���aҞ9kP�Tql���bs!V�v��L��f_�	ij�0�|��d�j����* ��N�����6u� Z�^�U
�ۜ�rg��ԡ�%�'�	�8�Gų�����&���.` K����H.���TR*9�[p��MLMá3�b��R�u��@���$~��N֧�ݽ��a��o;��]4s ����zCS���qw���<���v��_N3c%@_뾸�,�OD��b��<d�%|�Z�):T�v�p��<�߼\��B��>7����j�CP��{��� "q��Gԡ�������O�×b ��_G��Hj禞h<r�b��5W��7jj�3)� YasT�n'���[ ��T�$�7�H�J�`o)[N����2(=:�C��T �o�t�|�_vhµ�m��r�zL�_�It�����2YdL���kC\#&�l��9�lOm�*L����^ ��dr��@�6��nr�I]�a#��TJ�\̣���M�l���kn��v��}�O`?�n4�.Z�C�|�i���+���>th��� =���[���mFSa��m��b�ZEg\������"�*���� �F*�ڷo�$�t���ڛ|��7�d��������<"'7ݩvwQS9/��i�&H���7o>CH3�K笡s�|���Oc�\��ي�x�߈�n��SZ^�G��On;�I$��B�e��{`�}u@��+k����֣z�ia���-_�0�����D��8Gr0,�e�,NB�ի仱�z�1�:�?:::PrZ�*�҇o���;xh5 �Q,)K�c��y$�K��y��α����H �|���;i��=�֎8�<�u�\�>~7��r�:@a��Ī�Lt)<�+�x���~� -<E��� �R������byH�f�}��Y�|�C��I�xQ��Y�J���4�+�,i$����S
K���S�W��oa�⊣�j(�&#騸=���O+�6z�2�wbJJ$�!Ã�:`�� �H`۾�-����хpD	����1+�4�M�N���2O����u��g�`v!�.��).��ۚ,�>�>�`��򱱱�|7�V�$#K Gndr$Q���s7��b�r��x��i]*�Je7]I��E�x�w�I}�Wz�r:15�#)�M]�������13wF��p`=Г��3�i�R2J�1S�¿�Bר����3���B�u����y�o�P5'L⫂"��m���]�,��@]���0����چQȭ��m&�v���!U�!I�f��`%1ϛ�� �E,�wמ�c��WeK7�\{:vba��v �yq;{ج���?�li��c9�u'� ��7B�c�I=���Y�dO��������z��\s���I�Oʻ��?Z�K��(74����k��T�Qn>�}�Br�aXL6C�����|
&�3��s��;3��u�}2P���q":=��v�Q^V��KKK}���,g�H~>�Wu}b{�v�Um
zڷ�	= ���~łf�녮}ŉ�Q�[;L����Id�ʞ&�9?rNe��ɮ��zG ત$�)8�F.�K��R�LAO����3��h�ݦ���#ebH`�����"����8z��K��:���z�G{V&a��	XCG���3ؑ��Z�.�.�4˱�è+��0��M��������v..j���ٓ/K�MU�}S5�[1_���+�W�#����%K�C;OD֘�#���m��0P��]���!��a�D�m��;�`�ı^8�T�¼,B�}=��T䕖����S;�r����

_����\�F�x�� �Db��-�h��ύ�&�/�{*��O'w��+�Qp�+��ܽkT'�!t6�57߆a�?�n�	zMM����)+<��s%��zx���{�0d�=���Ѹ�M�!QM:�+H�Z�����H�=B�l�ɧ���C1��Q3��*�>;Zjll�C��~��JA3�$�U�B�E��o�儭�#Z����x>_��aAg��+��5�<��c###K��T6�
iа�U�b���#����_}���s�OvO��)���>����)��Q��xC����B�PŹ��ԎLIS ���y�>���i��D	�P��/����t���Z�2b u.�mx+���Yl��ɰ����9��C�o{��.��
I��j��kj���<�Z�WQx2%\,�cm��h́���Ka]�jʽ��� 6}A���0�O�ݠ���UZ��[�B��=ox����vQd���� �W"P��h3�9@�%=�T�#����0C>���Ta�|�d��^j�M}�r���Y�9�899a��Ә��F�1�X
��`�,��,08j�e���PV*n	E�5;kh^��� ��U"�j�权�i�f�!;�)����d!TH_P3���<o[D ��r�-�F�FTH6泲��f�� �~�x�)d9h���9i���M-նe�ݓ�0c�9%�C[�b��~z<�9�3$��G����+��J�*��{XB����"<�hg����7��p�֜��yR�2"�,�� �u� |�`��y����j���g$�%LF�����3��T�RUZBf�U���l@^�����?�^2w���$tK]������T��5�������(Rهr��S���f��$�J|s�^�jtv '
º�x=�I���"�Vh���|~llj:�t[���X,�6=V�Óo8)�^8zKN��s�$u*��1�xE�:$�G}�A�nBЏy�ׯ_o6ʵ�ʗ����#������̊1��caX�"K���̈�4���n�=vl�}Kjtfff�A�I֞bW���X4��c�[#r7 \C�V\�,A��XZ�,��Lj��
Z덠��ĭ��{���8:2���y�b&�8�r��_ϣ�t�� C��ya��Q����6|�y�Z��h�ژ�J�j�E�@X!Ơ�<&�~��VӜ|*Vc����V�^� �Q�YN�·cV&O^�P��~�s���IY4�?[؊��h_��v|�'ߍ�,:-�m�oIݐ8ӴY?:�20 ���fC�7��ֆo��+e�`��ڮ'+y)M����T�
����/n�S�x�x��	u�s�E7��+�o�)sH���!�����9tfu~�C�����$x�fc����jV|�ba��M���5����I7��9�4�� s:I���C�S�rH�N�ޖ��o߾��"K}E�\^�>Q$t�v��f���b�(�~-���;]}A+e���0��KE��*r�:��y/�]}J���R�2��6k(����������L���R���v������dȰ���w��[�l��z���R�.E��)���o6,���a9,��7��B$@���S�uN�eW�5Fqq[Щ��W����� #�\�<����^��ȅ_�Nf�*�z&����8j߬�ډO�*Bf )}c���˧T���`�4����XaKٱe�"���J�����8�R���oR������;�p�	��)�mԕ�L|͗����M��������n�p1���-F��s�[w=���([x�5�O'F">>~�s&��B�2���5��F����GPS��AW|��C�&[�Ғ��1�� ��QdmAA:�U35��4�`�Mi�v!�`�m�t:=̙����B�oN�W���A6��5P2��W��7��ʨ�8�J)	�7��qO48I�?T�6�Ec�hcc����G4��XDh�UB'�h+�3��ERw%FW�?# :p��e��
l���VM��;dGd���i\���"�����BM�!��<�ui�4�s5���H茀'p3���j@;��$�_44��y<L���cͻ�I�<ͫ��]zْ� �D:ج��n���P�����<#�V�L��y�V���q��?ʓ��v���]Ͳ x;x��bL:O�4�=��Q��crr�3tS�n߮E��$h�Tx�q��?���ؒ(>�	�HRH/o2�c~��@v�T�4oA���H\'���^	��!�]H����CbKx��4x�si� �N� & ���W��6� Fwz�����ox!�&F�!�BO;�8��: mU��7Qh=Fʖ��H&#�����P�Ԍt������1�W���V�$���|��s(YX���ί"cf*��5t/h7:x���E䅈�16�.#�S���A-̙^J�>���Lf9%�=Üa袣��>�45Q*�(:�g/QW��0q _��M(P[`�1�����
7�hr'�Zy1ncq�}���N�u�OCCZ@�� '9����^�ɕR�Ţ���5��+S�'�ƁS-�4��ҭ�b��9���IJ�7_Ns ��_����.�Bi׉e̡�)֪���f�y�&���^�L�@(�̃�e#[��P�fr��	��"y b�k�f�_��eY����嘬��
�Z�4N%�������M�����m��vq�CZ�7z�,��I ԠS��Lt�-f'qH�*�ů%ڕ��~���UC;��G;�z���9�rj@�rf_8�= �f�G���A�Xc�<𨁽��ކɛ�/l֋��ފ�f�?��&gp�ig+�\9P:1hah�5;�=��a�#"kdFŇ<u6���J���&S�SBvb����/�XRv$%�,��ma����5@O��������\4̥��Kۙ�T3h��9]]o��E!o�d�-���"J�W����8����s��nʽǏK0�@#/��S(mIc��)�=M�7<��;��M���>��mz��P��?JI�RZ=�����h�H�N%7~=e���J]�UR��ۮ�V|Sq�3�T -C]�_s/��`�����o~K��ޮ�d��F�2y��b�*_ϛ@TNp��T|g���t��>0�a��ѶPK4F����O�@�%P˩�u��ϼ�Yӳ��~j��fP�~#h�5O)�A�T���n����i��}�YUt\\,��S��U-6D^���Q�8�9l�'�zQ�����h��0����l�/�a���|��R!�E:w�k�I�$���p���K��ߨ�	^�[����"�^t�O��nQ�:�B�A�!��+A:��)�Q�a��&;Í}���%��Qp�����&�B��;w_Z�0p#�7h���1���[$P?zb�$�X��k��5��e�sO�˥�2�`wQ_;O0������GS(�a<�t=ЍX�ޖ�b��c`e�)
<2�c�s�}�����Хu���o�ai�2Yq3��n�T�k���x_9��ߑ��]�Yn
� ܔtceF��w�=���M�͵��HZ��1�_��"]�V��KA��"P��,�^u����T����p.�*��$�S��St߽O2���K(�| ����u�@�I�����r�ѫS���HA�V��~zQ���C�Gmm�������^}�x-�8'��\�A{���z��۠�pG^���K�7�>|�l|����q�X�k�pE���*7w��5��&���d)�7�P�P��*�P1�M|����Fݘ��XR��j�z��9x�L��H�m�͈��sH�E�֠�"?5A.�r���̲�O^����04����c�S=E�x/p�D"t��vO���)�^�x��?��!څ�����wM$) K�q���ec&�����!��E^5;�����ҫ����?�t��B�o�������]�x�)2%��/64 ���3e|�	���A�����z1ϛ�GC�����##.=��G�����/b\{y�,?�`�\�,ggϰ���@����՗24׶��~K�s3���c�-��Ik�=XU����JMЬ3�B뻌���8��P�v�-w��<��]	�Ç)�Og�^8$�.�t�-�Q(*.��G��-����L�R�(NC���Z{{}9=I�����A;v�D����������s�J�/_�~�����h�J8��)?� ���������@��X'�W{������]��H]��`*�`�w;g���ƌ�/꿬����I��m�蔾������ݻ���-BL-p������X;5u�իW�����6u��F�Tȁ��pHe���
��D�B4��j�p����P�H瞲��ȪJ7���%��_�-/-�$�3E��"�* ̹��\geŶ�2S	t;���`l��7Ͻs�s�:Q5�q��-@��K��X�bYK���9vnmoo m?+˹�9�K�ڍ��bK�� V��s2V!1yD&�c�>�k]�N��5�x���ɬX�R^1�Z�F�������Zu�Q:3�	���^�~��T�nW!ڐ
�\���'�G6˹	��+�Zs3jg~�����[����+�͘܅�n<g61�6ta	��$����ccو�����.SB�p�!����:�ؐG ����h�L�S�W�����ܻwr+�30қ�lش3g��Q�o��H���B�~�7��hȏ@g��gdr�uO����h�kE�Q�+&t/���##�%~l�a�-X��e�*��6 ϰi3�Νhra�N����Wхc�>%wz�3�{�-�D`��jM�A�D��!�=�GBSD�%ٻI
�5��#����U�%��ڧ�*��]��#� I��� �%��Ӽ֧�A&i������Wβ���Y�>6�8�T�wuإ�s��?�l����>�D���ߛ�9��׎<a�Q��M�_����p;����۽��?;�(⢏�,ge�rTC�d�2�� ��*��꛷�p���sO/{~?���?"|��X4z3�ہ�
����m>3����?_�ϊ�yV��ܝ
.W����ꔃ)���:K���!e��Ȱ�Txw��^8̏ѹ�H�� &�<��c��D�B��I�J����Q@@��H)w�������X�EC��Œow��P��!�RjJ98[�n�Δ���П;�a���s�8~�:]��f�I�"�8�NH��ҝvr���BX^���� ֣����
�C�������j�E�tg~�G;ٞ62㐸$�������6H�v#]�82�)#�5Ac����Չꛎ���zE#���`4�"��(�`~��{I3��L�����~�ey.�{������-��7�m�\rڄ<).�G{Z�M�t#�k2�O�������eLUnWK�R]i�����MU�$ü��v��BS�ΝIݝ�S�᷿ߕstu�SpQ	&s2�]�^��s]z2�x�9sje�A��=���Mr�M�IB��M������
�.|�r�K}`+�S	=c��b^{�\����>|J�8tW$�GsP���Fv��z؍�]>�6�ٱ�ŧy1p�S3���K\�'.	�L��+GZ�ǣ�omTA���@�u+4͆�k�?�4Ìv	Y��j�/6 %���-#��|���J�}��V#l��R"����wd��[�{z�tzΔJ�b���
��{+H���c�9������^'�\��ܾ��QϤ,7�aC�]2w�N�';��/>B�Z�E�h_�N�w`Wa��NN+R��������E�'~ExSY���D8�� ���V���3�6ю�I)\�2��UA��?i{����	�m���6�^`��o��In�n��Qx���uQ�:��D����F�k��Đ�נ媓(tSe�'P���t��y/3��ր&@�(�;�_>��/�rrr"֗|��رa�����W�̋��{�tKWBRR�c�O���{n���9����V��PwO�U��;7�;�r^me�����ߏk�/�<��`����$�#|x�tc�u|<g���N��d�MJ�AȞ�	@-GN�����)� �pa�2t�_�^��"��'�,C��r�c��r���P���1UN)����u�^���\]�b?��("��]�hq4�B1���V��)�|V/p1��7�qP��Ι(~/��3��G��&�!frYJ5gn
d�;�6$��#�--U&$G�T���ff�f��K�B�EEF�U�l��~Kkt^�z��"��a�ֳ�i��Җ�4c%�Y.|���3ߧ(����Q�/}2��F;��:�\��
7z)��q�v]���?f���ţm���q��X\?������t��'�Vm��5l79�R��e���M��|z�&z��)��+����>S3/�1�Y�?&��R����gc�����,/X'ly�����f�#`yϮ[v�&��Fi��X�f@>B=��u;"��I�CP�I&s'0*��Qo�:ۙ����:2���^B��@*\��q���O�+���pn�F�W��
q�_��閗���**&f�U��Q����z�ZJ39�K�Ts�\`N�xȹ����b'���I�����LL�@ЪƓ�����2~���H���ZVU�BȎ3x��Hj���p���<C}3�X�E���ˢ��<cI+�K��D��6������i�;���ߚH�Q��ke�u����O8
*xX���	��cޅEEOu3�D�[G@նB3���޾�i�0�6d���
��+UyP�@u�D����'K"�N�O���U�i��	.7@IE�V����O�f�|��Q������!c.��5�1h�Es����$1v���Hl�e${�F�Yvq곲,T��d^*��vU)=镏�o�N�%�V	L�d2��# ��W����Q�τ� �i�>~�W:�����3�1�Q"�2W}���h.��Q:����ë?�%KiM��u/[����-[�Eƞ+�"E0�*W����B%��3Ϯ�KoIN���g(��t����?x���t�N\H$�m�Y8�Zdg5��q�\�^6=�_����XwL�C%Oǜ�s�rsp�Y�b?�8d	=QZx0���)���j8��/�~q�Ι���͢p���(�#k����W�*�Pt��v)��0>��Z�^�r,Bn��=(��=�_Rx����&��_1q
Ӊ	��T7Z��aip*q�t$���rv�0�砂}>�lX�����?.Y-.�H����z�'�B�	���Urhׯ��i�t�A�l�`Gw�?�꯶��I���V��'C*~я�Ȩ����?�qk�>�c���ۓ���l�5�D����������H�j���-��S�5�Y|�|�)�1�/�ʸ���o$���!��l�J�Y�_��M:WEW3���58yV4�X�q��������@4��3`O�`�׀P������� �
:12�-��5�:ѕ����)K]�;�k��!7_�ۤ-��k�˗uLx��U��u�^�;��ļ���d�)9v�=~�0�i��/_2퍝��M���g#x��(��4tc��f�u�F񈴽mD�v�gm�[Q��}��7���`�s�5(�LG89�?5��U��N������acɢ��k�[2]�i��PU�|G؆2"k?�,s\\��/���j)�Y��B���9����P�#U8����G���J7h���#��1 1�n�Ю�H%�Ĥ���!���ѡ7�dj�<p��J�Z;�s�qo��tb���i��_Me�/���e�ݔ�D��������+�h�Q"��T�i"I�IY^��_Ey�:3`��xD���T`NpU�ڑ9�[���̘虱�)T"�#a��k}�[b%�2<���{���`hVX��?|	��-�kO�&S�{�;S���~Vԍ�QMh�BT�̠8�X�g�G7��vVcmFj,i8 L�3p�	{�x~fpvq/n�ߤ�Z�z@HH��K�{���#3� ͏��k�{N�bA��S:mxbq�An1ɻ��)�αTV�.}�xU�*�l;��^�{�	�Z�ݱ�H�|䖛Q��Z��*���;��y�LJ�a|p�X�cEs��L�i�9�Q�֓�>�֚�}F�wtgH�[�!&ּ:s[�s+�_A����n�O	����Pȭ�d�����~��ʅ�OG�;�L��A�ڙ�`���_j|o^T\|Q�6�a��W�H���o�2����ATO!��5rg�)1�/?L��ib���z��k-�9��Kh>�	��&��Q��w���P��#���Yo���W�������RVl����Vh�X-�4���q�+ב��A��N/g-�mpz�5>]9r�>�F��i�M6PSxI����a��y��DED~�E2�s�a��Nc=�~�		<RWٲR3R%>���d���\�MD+ʾ�u2��$j暛�knް+x�%?Y�!1�����6;�q��c���w�T�gDl"
:��9KNMg�+4p.B<ƑiM���ͥ2w��UL��?Q8t#�_����*����6���!�����U�u����z�Դ�y�pAI��ݝb1s��Y{#W�4*�	�zjiXƏ�� l���)��e��az�˯��*8;��$m}XA�0�����*2)�!-�$.eF��q���L-|���wo�h�Y���%��A����&��\�]��í���t>1_���_^�ˍLL�������Pfo���/!&ځ&���D�����(1*��f���ڕЂK�x�U��G��3�q��o�	Pu02�ӗ�B���G����DFOs3s,,342�h���\�P�q;v{t��ه�j����]~HNh�+������^��G��`0��E��G*)��绰8�k�j�o����vI������qP�'�����䐩&D�e���37��By�L��@��ԙB�B{ky�����]��0�"qkB��[/3X�]�-T1����m�**���?�)B�m�l ⫟Q@no'�:��y^���rv�(Y���"���h�o���05�r<A|$ݨ�T����4������2���Y�mA�\z{��D�Aߏ��d���ޮ}����R��n�7U@C��� p��Z<��GF[5'3���k9@���L�R��Wa�������5g�N�����u�۪�6��gƚ�
FNW�&C��|[||l�V���L�np�G.y�V*�d _��Hx�g[ak�p:C��UNь�;!��/vrқ�_ p��8��`%T=�{u.xI�7�͕�͠CSf�V(�*�
�I��;��@~5)�V��ΌWg�Ţ�;"�;6�1�P}����P�3�o�}�^6I�1 �,��p�T�m�޼��Ј��� ψ���͔s{+9
u?Pl��L��8k��&.D���z3Q�w�3���j�3��N���64�scn�������j�Uq@v�U"c.-n�FX����+���}k}$�+�q`�\]�ſ��q��)ux�dT���}�D&�x*��+�w��^"{�����"���$�y1���)�e��|,�5C��l� ��_�{Ї==Y��x[ۈՇ)���z��|���#0F��٨6<P�ۗa��J�-`6�ҭc$BbH�YC�9��VV��o�wc�x,�,������O�9N�G.��m�꜇��G�ޫ|��� ~�� ��]�~�����7���k��������Ti�s�b�E��	��g�����H|h��IM��j��+��#�mޠ^���&��sb��+V��$"�R�uw}�O��X��+wwu�{��+��ۥ�H�~��.�]ۏZ���99�ҍ��s'�t�:�XR�|Bn�H�?(�f{{�����aJ4X��\�m�Y����Y�T�򾧟�֔j@�
é�Y�u®ً�ń������Qr~�����	n��Dl8s
�ܔ�EF���X%�f$����͹W�ޣu �촥Д �r,�P��!���^SKsprhs���9�JV�	���E��/�w��|��o�>�����	ݼ��§͋W�8�$��k>���!�]DJkw����z�a�۫�˦�M>h�?B$��6S8�	�TyV��G	��ߗ*�����J��o�`�zD�5��@���zb(�+φ=�}������G][�T�{�uM��N�@!{�F�׍a��99�����z_�^�g�rή���qx��K;ِ?z��emܥ�yU`hha$891�;�7T������"u�b�Sл4��mV��@/�%tE�[��]Z;B(��^�����_Gw�Ә��������e<��.U?ې[�靀2�ҳ��$m��,��p�o@��q\g,�U�q����l��,�e�]���ЃR���ǯ��?8c�$�Tq�_yU|6b��K���4"&�S<d��s']��9I��{a�mxA��u(��t�3�IVu�Wb�/Mm8c �dw6���/[��A�o�\����1i8$vZ	���T�r�[��j�,h�|Y!ˏ��Mꄡŷ(�N��L6�J��/�T���s*G�Q;@0 @Kj��o%��x@�Yz�	�����}-lu�]b�Ui�[��Gaq�w�H����љ�%�lH8ʶ�OrPJ�p��x	�6�|�:�4��8�!��zkڧJIq�:�r��'TT�q����f�a0��ݏ��8۫{u�lv�2��i/Oz,=�������T���Ф{|�%�z� �j���nVk�cն_��~&�ދ����l��W�[ �)���4�1��V��6��Y��)�k�r���3��-"��|R_����aa~,�7)�	�Ώ��m�I��#��v��I.p�ĉ�]�S@��kmZ!��?g��ӹ���^F��,����]��uRJ*&��(?K/i\�3H�#��M�u�_�EK�ZG�p�HÞ��Ƭ�Lf��s���B8��_x�NH(lSpo��0���o��be�!������Ew��֛fi�O><�\�J(�㶷�z��.��+��8�!Cdu�.��&��ۮ�G%�=�m>6+}4�B��.��R{�C��
�:�$G�/8�dw���&���~a��^���]���\�ȝ�j[�7��Y�O\��@�/f?���lk��m��}�3y1m4�SH�X�Ԡ�ڮ ����MQ�����+.��3��:�A�I�[�W��>�󭤆~���3T]G��Y/\��]�w��^s:����iOq��Ch���^���w��O�4�S:��x�k�~l�?�
T�'4
�>�|�Y��7-�!��q��\�8ipN����Us�m�c&��ܺ ccc�!!zt�;S��na6��-N�7���3(�U��>g�jao��1>�����r!�fuɟ..�U^=�k�/�s����|���G\6�?����W��ЇuC�#R��G|�-	��S.�/�*��Sl,\���1\�d���"&O��>�F>����[�5���ĕ������==���$�;�4�7}K�k�^�P�NP�)�b���$~�n�͐C��}Ƞnۓ��o m��|��jϭ��#k��gf��XK�г���|稤5Xy���'��kg��6�9�E|��*�#�:}�(5���U�YG��W3��+��nޚ�˝�!p���1z��
#��jj" a���S�f$O�̩����$�Z��&B?ޖL�>��6�Ρ1��<��k>�J���E�2h�p�@�1��� ��'���mU.�e�Y�A��ۛ*���J7��$@m���DCcm��>K[]\�q-��p)� Mv��B#�0VCY��j���S�Q��5�lIrv�H�K7�ןݾ�G*'�-~㙣H���\���z�:>�f�Gn,*[-�����z�K�YR�j>U���y0��t̷+Lp���?6o��ٮ�uUQ�܎���MiG�!�1u��ſ%��Vt|�x/��6��ݕ[��,XGE<李EO�E����/���_T�S�'[��������?��b��j��i����꼫]���WK��,�z�tds�O���ѥ%J�y��lՐ��9�I�<�R<��\WG/�8�z������Yͥ��&�EUà]��^'F�����T4��6i`�@�y��NO��w��.�{dš��>���&/�����"
�����o^�cX���;���&6����\IA��q�O}�%�CW��<��O�i�-��t���͐���2��B����;����7��VPGA��ڈ`T�`1"��A�����Ju�t+̈!��!E�AJ$JҤ�B��|?����u��de�˓g�g��>{�s��O�r8C]]ʮ�bRB�깡��ῒxju}	Q�y�v��b8f�������g�����Bj'�'`�ď�4*o�J�z�Y� ��k>����\���w�i�VVT�}m�_�Կ��������N���H���zK��dݘq�?������̄=~^���O&R�@Җ�	�Z���4��5*�m?d��`!�)��<xw����A�Zn9�Wk�rKl\N��ݵ�%s��T�U� �ݒ7O�'�x�Q(R��!~	��6[q��R���~������ ��q��m@�F%b�C��"�>y�x�n�ҫ�tl2��ϙ�� FN���i���,~T��U��e������ߞz����Q�8��E|Ɖ:x8�" �h��:�I4����X�UV?���b��ҡ��X����g�r�������g�M�i"6��6�a��7�G�S>�>Žc�P�w�ι��r�+�/���pE�����C�����+��8شc%�Ĥ�Aȋ��f�M ��S�+_��^�2���KQˇ�"�yp�j��Ɍ�d�({E�ZˇF���-)��C�r~Or���]v��
�+l���FVq�&��\�/�8R�;�Ԍ�p��rB�"�=�_�խ�)KWX���B�N寅t���W ��Rp~�5�(~v�ο�4�X/~�Yu1qI�'�F2��$cd@��)Z�^0h'_e��ysGҖ+�ޢWazf���q�����++��F_,N��#In8�&��}O7H��J��#��=*�ͯ����Љ�2d�������$��~��NP�DR�k/9y������[,&���$+9�K�d�xV���aYWU���7?vA���։��|�`������m��Q�J��(�%�n���Uv�Ck�i���1u��Q&�w��>�(�Y�ē=22��,�y��zE����@�az�
ӗ֌_*�N�#/+��1����=A�?�������)�F�  }�yW`5�����7c����ٸ)�p����X���������ū����7 8���,�����7ъVnٹimSp��*Bȍ��۱�G��J�g�d4w�f��f���(ﴃ��"��@ 9{[���8y��f�/v��tCQG��B���j�Ҋi�	�:�
M��ϰ�q�ħ.�Q��,��e�{��
�J��u?�L{`��-(��*�1)��ҧ\��$+�� �J��Z�5Oe�*5 �)��p�
�.�8{҈�!X�J���8��b�%���P(^��?/�]h!EC���H�UͿ��T���]�@�d����t��?��7�8��BFX�z��)����m\r��� �dL���I0w7����A�HUA�eV4u^-���!��`�Bk� ����U:6.�m ��K B�d�mB���,&�-��A�9^��;���o�1?6����
k��:��_Y(It�!K�&��@�p���d��uÃф��Θ!e��H�	�G��ς�ZQsk�����%�C��N�˻�:$ѳ����
��w��F� �� @�F�R�<N�cF������Q}�,
<��w�@�$��SE��
H�F̃n?����ߚ7�0lp���c���-	��f��,�R���/A>״��������6�����0-�M
<���]��T<L��e}��s��4����俗�� ���a0굍q����u�e����)�+��/�� ��R� �+^��U�����ߥ��
��}_���(`8��e�`� A��t{�P�����f���!"�d$�z��#P�]EV��%�9H�EUz�pӁI3h4Ȓ�f�$jf􏏏?�J�A�b�Q�F�9�uG�\��.��"��H~�։# E���ws,�-����u���w~�	,�����1���l�-埥�}si�-�m�������0�-���A�h�%�P���h��;Y��#5�֣,��\��	`!��~��G!E_>K��O:� ��ew�nGW<�'"�t��Hdu�D�p2o ��F����]�.�� >(I2(��dl��j��Au�wVՈ^�Q�m ��������ʎ�:CZ�,�ͥ���\w�3����� ����9�@/�ZrabtDjU;���8G �{��$¼�4�;w$Q��0�K�oP{>!�!k������	���Q�M_o%Q�뭴�n�+nuY�@���-���Af�VEE�n� �TE"(,N����J��f�UR��;|e��!��bEÚܵ&�$�e���D�~4 ��dF��`��&jNd��1MT�6��:�!g�e�M�Z�f䡽ԅ�~��Wf�s�%KV�^��]��ݘ���+��9�_����ƹ�Y[�;Eod�d�-��e���q!=�	��ȷ���:/|�l����Q�`���D�MV����3��W�#�fe��D�g��S�h�`�N<F26}�yz����G)��dD��[9I�U}��%%%`є�H>�#`߆�VF �2x��൲ׯC�Z���yvDYE��"b���Z1��y3*��]T��n�Jj���qR����ZW��*�b�˪u��M��s�ٷ��6P��F���WA�Zn��1�7+Q��G�Y|���B��iI���Ew8�G<�.>T||n��g�?�>������J���y����H�Y?�˺��i:q5��k5�#ȆF�ז���}_������9�\�!!�0�k����Ю�HO6���g+{خ��F[���猪�#�������{�u��K��������QUo0�A�R��ؑݻw{��@t[��N���s��3�֡��w��2��2Լ\u����p\RtY��[W��F�M� ���nj1�ܔ��w�Fg�v�Ai�~�֚�#��h�)pzF��D��Y�t{�+��k/�j$}�%(Iw�[�~&qX�{�Jl:`�]IlW�ߞ�����@��̈�.?ᅗ��<&�#������>9ɮ!6	K���pT�)@�Ź)�����@��޺×���ȵ9���d�-�qj>ӄ�ϐ̬A ZK�����g��@��?��O�#N��3��neHt����}�K���׏B���$P<ӧ�{����,Ev�m�3a_�}���z��v���98{�w+���Ht���Zc��F�S��P�(@��0jT?Y��x�$M�����I)8��0�H�آ��Z���ĥ��>�X�Q~���ē U|�<��:��G�O����>A�������}�A�}���5��3�^��-�w�<]�bʜ��RZ/+�I���=�/�jż�V�*z$�v�G9��f@Q/]E�!�_9T�:1�[��=�U�g���-�3�M���ǟ�Aj}��G�����>$���?��,e,�L�� s)����$yb$��Z۴'�������"�J+�,w/�lb˩4h<�����4�3?�����A`�Q� ���*���9�\|"����\ 	!����Q�ɸ%op�M�>�X�]�ԛ)ZZ>���6�V�ҩ��[;��1��	�gAY`�h)���ڥ&0�ϣTY����܊
ڲ���]�O?׳�cIgh��s��>�vfa��,��c��yg��"I8��>['��T�~��T�.
�T��8�I��͇e�E��u z�Y��ݐ�ġ�m���|'�
�kbd�A�tz���$X;���_��@�:���;���ӸUrx���"2�:��O>���# y]��{�
�f��\�}DMf|�&~���z,`���u9�����<j:!�5��K���9 �X$�����⑕���?������}�|z�j���\ZÈ�6�$H���g�P�qv���'^N�K�~"A��(�ϑke.;|�����C�#�������d�Ê�! ��.�����~�W�]�d��	:{�[Q_��Z���b��+U�Ϟ.6��.c�
Q��7ܬ�>r�jއ��ˉL}�g��,�7�p��*�ɀ#�[8�xH��}IFyon��M޴+�zk廍w���ξ���_�,J�BK %���섾�`�q���lɆS��YXu^�I�kL��'vd_e�1���GC��Qr&��@���o���̓�a��$&P��L���0���LNN������}V��5c����/��ڋ%�2��6���G��Րj�.x�G�c/�ս�8��0��_��8"񘌚�x��k��6QD�z�qR�����Ꚛ���oQ+�a�:[��40��6��a�>�u}i�}��`�(�\q+1I}8 #��j�NuA^��ێ���݇�?�]w�Դ���֧����Iޟ۸�d;$�2�%?n��Ã�@����;�ۻ�W�f\8�&���k�&T�1@�j�D��c���k�$�O�8�'������	C �H]#���ߍċP���D&��� [gk��m�ȈNa!ǝ�T+����h���^�٢�F���\)_�zw��:O � �jx���<�niI��OL\Zٟk#g��:E@��Ja*$�s���H��2'@�	m�-����%�Di�c.DV�y��L��f,²���X�f2��0����K�Ǐ���2�������ك�+/�?Ǧ�3��*�-H�1�,�-X�(oB��1���0v����u���`��j����kpDxxڅ�Ja��N�W��|.^�s�U��ԙ�I��dm�Z`[�����ط��U��"ӻ���']UrU�ML8��n��7ͧ�����]0��?�V�WGf��g��͝�ԒY�ل�!�����b ��D��L�K���!�n~�C�}�8�l�8�gΎ#d��ޅ# M()+�����˫}���r*nu��p�U ��z��g��Y�Y����Ӌ�)bEe�":�
uk�=$�=�Hd3~��W� ��4��P��GN�ED�NW��7�ǩ�U<	�������#���u�;�Gq�j���l8�^��n���4a�7�;�~k9I���F�h6u�pp�i]��u�y�39lƄ{�H���nؗ��"���ܟ����`�1D~��G��#q�HksI�}]��3PAX�C�ѡ굆4�ӟ1.�)�W���<�i��NN职:�*M�����3��+��.ɍ�9�w/<���S��6�U��"�����u@;}�	/�������	p&��{����]���2���[��G����bP�G���2�{[�����/3����?��ӃhSki�ㅬ�[��ܼ���>�Wk���V�?D:V�u��s���ݸ�� �V��5.�a�q�j����'�p*NL�dG`�9��0D�s#�u׌k��^�_l��Pd��UL�ƛ33a��ᣥ���3���{{��Ig��&/�zEi��]�7k����"�1õl�f7{��O#r<T�rz��ʕ�����0�z*ֶ�*�'�-BM���u�q}�����ټ�0�@�-)�LV|�a����	L�X�s����oe����4[��s����Aov�S#M{b��c����v)���:��0̞y��[\wM�$�5!\���<�QK�b *�2�%�3f��¶�f�z������bj`]�%�E�\$�n�����#�R��n1��� Ѯ���mq��9#��z �<R���V�a"�\�;_�ߔ�-	!]�j��!��ԫ�}���{��'L5��?�1���Ev��VF^8�^�2��+�\a�	C7�ٗl�cT��\Yk���6?B	�2cц|nf��["�
�u�!�c����c��M�%h���OR0����2�hJn���]sA*�﮹QT9����J�.�rF����o��B�7�n��VDTe��Yԕ�]3	\���	+���CSʠS�����g�p�Z`�k.�&�c&����>��D�s�R�ʹ�U���\x�!|J�Yr���{��"�s]3T[��{W��G��;Iv�n�-�Z0���BVe,�ZA�g��K儚��!L��U��'���l"U�Q�`�$7 /k��m��:\�Q�a\_	c��[�2��,���
��{~sl'	�NĪ|�n�$��"R���R�YفT96y�1��L��c\�O^�f`�a�{t'Zź���w�W=�B�������0"Ùb��W)����NDF:�&�Y9�{j&�8���:��j3i��O��g�h�W��:��R�Y-��T�e�
�j�Y_�5yY6�z�j�����<����h�F��Gp�uj�pMÏ�����ܑ�D�� ��hka�B�l&��b��]L����V���Ϥ`+3{G��]��-{yxhTd
Er����"\\�[��b�z&x�Ӏ��%� �d����׌���6�������P,o��Bp�7����n�ָͤ=i����X�Ǽ��1~(zt�(�SƈL��B��:��6��[�g#Xmq���DI�T��Iʈ^%�Y�}l�cH
 �񳙰�����g;�J�L�-�^"�����Ԏ]ų�=�T\G��wAQe��!O!8�
�S`��������ͷO(W�M0��Rnogg�p��t 6�'$�8w�=6� M 8�ʁ:j�ʪ44����(]F������Ʊy8�q��f�<I�-jD�&Q����俟4iT�|��~���������X*�D��W���N=&�T8��čj����Ij��$�I.�\&�Lr��2�e��$��/�.�C N�f��_&�Lr��2�e��WI
ٍ�N���;�qC�Fn���7��8�j*´��ҏ���T�?�~���������#���	.\&�Lp���gs�%S?�V!���I��<��Ҏ��Do�C�?�]r�r���'�k�Z��&�~4F�+��ѫ=��:��BM�L��4ū�P����$�0�Q��7K�:أ�-��#y����/>_�����rI�:�����j��Uc���e��UI�?U,����;�(��Q�=���÷셛=��D#,l�|a~��� PK   ���XhT���� ċ /   images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.png�|y\����Td�D�+!*ZD˴qk�J*E�B(�F��-��"d�V�j�s�!5hE�(��}�]gD��<�>�_�^��m���s��z_��u�3~�5�7od߈�`6��(��`60ƪ���/�싿��8����������7ت�s�`v�F��)�����vCQ�������/a��Z[:�_��$dcoE�a�`x0�
�u��}�R�8��w��`��&���`>�kq���x�i����-�S���q�A�rg1#u�]�u�\��ʖqѽ��D���A��뗬M�N�Wj��S�1N�0�����^a0-ⷥ�^2�;R���@�z����f����n��=S�u��x^����:v�5��+�5����;����w������;����w������< �M����R�̼��CwR_y��ح�|2��t���S���]o�[��}��C&-�Y�5�	Y|�F/	}<W�|i^u��b�ud�MK�e��W1�F�]����F�I�G������&Zꅽ��c������7����Ϳo�}����������lY���и�vKr������?���dfE-���aƪǛX�nd��z��"��&�99����]�ʎ>��4��u�8�O �d�%���	g�}��&U���x]a��{+�;;�٧xՏ������ZB�����A�ca投�B��䠏����d�������l�i
^�QHȤ�����[W����9�9�nj賍q����#I�_��Y�6l���xrR��Ӯݙ���\�/_�Ħ�:�|lB¾���FB�q%%r��~ۄ5�*����i;�)B���q`�~�*���;gF��:+�l<�'�%o�9�I�?�w$�+j)��˫�,ѺU;�_�vRU8������Z̕�~�!rMG bf(��ْen7�����^ &F��}��l���^
�ŚU����M����{���M�yWVRPPP2�9A-�s�[���4<��ʕ[����!ܚ�v�������lb��ˊ������x��e���fii�����C�{����ޘ�׷�u}xv�n��Z�iĔS���߄{ƣ��yL�Q�'L�9���\-q|���M�99G'�~�)��璛����Y6%-y�c0+� 6&C��uO��\v�zK�W��a���[k�L_���g����sRv��Ǒ<St�fF��d[h�J�l߯}Jv�OP^+5+KԺh�J�`{�����ʬh�}{��٤]&��oү[gnjʣ#�w�f(A�N��ŕe��>298##\Q�jtS}���$Q���7�|���	N�f���k�:9===���h<��uA"������o�aDј��\Y�v�
�U]�*�SSSsbb�≔C�An�U���vRڑ��k^�7ݺ�3���k:�H�WllB�ڔ�>8xnۏ?�{W���o߯Q1?\�=\<m�6���˽������^ϫݧf�^�L��@vp�4��p1���5�u%�m�B���뿼��/-�K۽����I1��$�]��WX�֐�J@���Z�;hTp+-�M\կ��r��Ü������~]�!I��0?��f���󱣃;��ACC,��������l��Us}ͳ	Q�J��`�mk�������\gF!�?77��au��[�I���%6��76oN�.?��֢e������b-��3��&'�sJ��{��p��;v�����R!ս����r�#̓㐣sRY!«
Φd����hur�����|r1�;�l���M�Qd:*��D"���rdY6g �&���^C6dQԪ�U0�h�i/�^
��]Anb�.��������?y�ĉ��Ϧ��Q��[��;^��\�Ӟ�,��_;:ǉ�w���>>"!Q�.B�+ڕ엘�H=қ�w6�t�,/X�	�}s����6Zǌw�ڔ/,--=OM�c���-����A���I�'z֐x�;�\&�KܜQ@R�.FL�Fʝ'�͇ۋ����b:R��Mi�;��)��L�� k���;'�MB��m������[@~�	FٽV�S1��Y��,�3���-	�'��j�Gf��ή��Q����RT`	l	�^�4�$i�]e@j/��~^��QQ�)�vLJFFF|I��.y~W�Ǹ��{�e��i�������335�M$J���6:]�,�4YZ�H���¿�n�E��SR���eV����T.f�}v�0�ݺ:C6��G!�Ĵn��p���Q%���uuuN��������/�Mca5�=}��o�G��~+!d7$��#��H��n��F(W��8l�d��G�V�8���.���˺֘�4����ݺZk:������Հ�q!r�,�"0����l����D����|�9MG�A_i���Q3Z�ɄP��������y=���7��[����㲑� ����Ӆ���c����m�/]�v��{�.��hW!H�g������O��:�8C�jr[a�XwM���=Z��;�vG�ef
���h�! F��-�a�� ���d5��0�!�sww�Y��ʺZ�x ��T�|-��KJJ[j/�.��h#��N8��JTfm�y�?��s�OԌ�%x6�Q�jn�'.[�TI�	�]o������ͩ'x/rߏA�-��6O�=�&�z�x��8_p����C;�ߣ��E�/���Us9V�ºH�o'��ЭoM}C��2�
m1Qd�c�b }��~�ª �	��'���-+>�����d#C[�j5)b�ޅ���e���G���V�E����mQ���7l狧v
��g�v?2b/�Ĺ�G&k�l�ׯݔ��dIOv(2!��jf����
�Ľ��h G_J��?��@ �h�Y�?�m��I�^[�{`|]�I1�ʻ��1�N^^Z���|���@E%%Y��j�^}��`q�����J �@��]8���fn�;N�'����������v��ф���1�@pnR"�6���O����z�Z	��<f��8���=�x#/���?~Fޑ�����8���f]�۠����SQ�v
s:��%E�%���tF�.\:���I��/�Ja���;[=r$ܥ��n[���n3ʱj�/�hhnN���Ɯ����oC!*~��A.��LG�[	h子2�����Q�uj1@F�!C�=���|�ܻ�.��5Y��\Z�c%�@o�:<\���	kD�<�/��ikk}'���o�!�v��% !��@)t@L`C���\��L�V~�X<�;�
V-�z�Ȇ[C.�?��4�Q��o4�p���-�Y�	6�cC3�V��M��� E��{ ��P���-¿��=�6�"�M4d-t�L,���jB��R����D�����Y�(	������$yp��+3=�<;�Oe����8�v�����Y��Gk7�!7�m�w��i6��D퀁/@�!��K�[�mpHyP��E�i��B����E�#�Kz'�nr��>���W7�?�]� >�������˓���F�f�LZڃRG��<W�~j���
2���]&�I\��^����E�x�g_L<�O����kF���k�a��?�4�z�y[��&�?��9ui��p�%'����uA;:Zͭ)K��Ϸ��C���X���NX>�P�D�:�bt�����#�~Jv�%�4�S �� �.r��^��B*��S?��!V&�|����(����2�b���kq��%�s����^q���T*?#jjj
t��O,�fVL3)�����F#��#�)�Q �Iѡ;��#a1{a�%b����J�|��q'���>���H	���Z�!R-[)_ʡG�e�����[�kܧ�X �թ-ɺ2�V��`������'e��i���=��c��f(��E(�W��sW=IZ��!x��g3�|��}^X(A϶�q����Uabj�*�(����4P��w������~Ϟ=kpeWt�?2ӭԮ��{��E��Ln�e��uD죭�(����KT�3����^:S)l�99)� �A�-�{��Π��?�í�կ��?~���Η=���CP��_�����"kFA|(��˿����dXN���m@��|j&��ʦt�8v�����r���&�?�OZ���lqn2�"��qf��r��n��v9��r�{F����wC��� F?*s'DN�z���H��_�����2L ��-RE�D ��m�	��8Pg�� �S�-�4�M�_�۾�
�7P�?V�p`rrr����"B�K��e� ��T�eg*#����l)�YR ƾ-h���U��c��xO�����uR	�8�|�KlT*�\�Fi�A,#U��@|"%&n�rυ�j�.�Ifs���qB�6��X��vC��#�X�n޼y��M�
���7W>���[%�l``@͘=fɣ�ň
Z��IW�l=A?v=0�V��?S�ɉ�
J��|TR'y��U4�jSG�JgV��ԹM�ʊ��/_��2����pE���p˳�ޮZ̈���{��1)գ��գR��FR[��r@F>I=�M�_�:ܧ���S���CC�ww��dX��WZ�Q�8�=C$\�� H9R�S�I�^i��U荌����39��s���`�d�Y]L..�����I���M9lkR�d�������(...`��)�CW��m�����{�߽��Χ�H�N�sǧ�N�0�);�:��^��V�WD�c��������!AduP����zR
Q����a���[y�z��sܫ�A�ժ�0(�I5?)�[��b�eA�X�#��G3-
>�����p&�rJ�o����%ub�$,��Uy9�=���c��׍ǚo�R���]�r�ލ��e��Ӎӭ�0^�/�+�,_7s��e���+X���NzN({2www'��5>e%X~4�d�ڵk���C���G�B�t�������r��囵tu#���x:5##��&2�nF�΃$�n�����R�	��;�ϯ�͢_([4�=�)uGT�D�5<��Y��2���=d�|��2�:�}�Qءgx۵�~�̽��h���ԟ��H�K�����⤻IZB�8y���PEP�c4 Y�N�g���i�j88�E]��9�r�I�]��e�Ϊ撩�Y������婎��ojj��ۘ�lIK�Dw�w���9�&T�,��))0��v�z�j�}͡?W!=\$���57�ܺ<�,��z����	���� �����Xj�F�F��_-����h#���'X�s�,�E֋�-��I?�#  (��Ǔ,�q�9^�֔��/$R��4� ��?6>�*=[�8��&hib�Gxx:��O���M�/�zӭU1��ꇧձ���7d����|�� �`0ã���|ڹl3�֌T����sM���#�&Ï�HK�����T�>���Jܺtqj�آ��G^Jj**��[o�z��y໧�؜r�E���x�!�������\*�XGF����u�A����6QS<�#�w�S}[H�/��YlBn̤�^2$S���B��C)��1I�d*�f-"��ɕ*�nn�<d�S;I�G�W��?��C���z׉�2٨Zl1UϏ�y�˖���HJdu��1�~�rJJ������e0}ю�j�s-�v憾��ٚ�0=���iC5�c��s�bލD��"R^Ϻ{�l�a�S�e��ZFFm�yTO~sdnU0�������0/�����}���v]ASs�y+
�<ON�O��n��0�l�}�Νb�Z9B��x�����H�#�g����S2��5�Ɋ��v?r��*��6�5��7�]m�率�(R
���I��^�"��L����##Y$ڝ�mLVOS0^4Wj-��n�M6*8���k$�7�<5Wz�D*[/�q�n�2�87Ox��S�i2�3�"DFFVs��	���N����d�#y�����kը4�H�f抗�j�f������v��z�M�T�aU8�i����2.:j�*�Q�q�}���r�s������Ʈ�m�����3�v���3�]qBT�,���u�������we�_,3��r��ܦ�ӭ�R�Q�sb\�9"���y���Hj0��jL�3�pv&�\��*aݚ`L�%^�M��Ή:�}p!�cl�K?�K��z���s��݊�á����J����P}��{0���ȸ�UR�ŷ�o���p5���T�?xP������s�[ �	2��u�̦zXdm�e]n����S{� x?�Qov!��2�|QؒD��"����A,
�I�cJvuR?@P^�o�娭0?�(.���������Q�˟�7�
O�QM�A�Ņ0���  rST�:�<̿�8����:��CWW�e��ݟ��+�;�N�ZGRx��E!I���f1�����8��Dq"!����[~�U�$lb'�@�G����d�E�����6R������pȆ�|n=]BWH%�T�3�i������c�+_~�B6z�T�Unn��p����!2B���7m"z<�����s����!������{8��B����qo�06����ʹ_3:������'r�Xt���39��������*���,����o8:�؟8~�833��ww+���1oxsO�03��(�K�����'����E�s�.�aY�DJ���0v���q���R�Xk:���E��
����Z�0���>��uuu!O�x���C�^~����CA�]��@0�c�Ν;�&���{<�<D�@�7g�̰�9b�ޠ��q����!��͂����Ό�����h���w�bcy�N=���4�y0h�|�8a/�&�]a�:g�N�g�Йhkk��r�좙�,������i�����A�a|��a�����5�[g~?�OmvCfLsYqA�;s���G>;q�����]߇g��DB"���%���k+t����(]�t�T���Ј��xUp�m�\�E�g�'6������.��/�X==�Wyyʎ�ӟ{ݿ���d;� )���l-f�>+�����7����&1��l����x䞟g'�$2��0*��߆ey./��zz��%:�EǸپ�������,-���{aK�"M<f?��Q>��+IL����\�_SIM��s��21I3&���	�5�k0�]�}��Μ��l�UU	�g����($QV�V���rc�D���e"� ���C~ʒ��9�����)�&9En㘟��>?U	����8�:Ɇ}��Ri��Rdew��.�ˈU��n��e`����R�0_	����x"ɴ?�|��W/�����D���?��������uH�x3�\�qDD�����d ��$��pH�Kٍ^����ۇK歁1I��ޯ�v],K�}��+W|��� ��4���R����"��=��T�/�c��JKw�,u�tR��x�= lX����:�S���qpp@���o���!������C������B��0>u���OK�`����g����CȻo[{l6646Vf��{H��<�����{xc�	gE�K`u�_z�B�i���� �:!�Q����W`�3�ی���K	�pهG��A�K����yB��dŞǸ�?׊CA8��:��y�����If�ux-==0��X?�Ą�}��c�g��j9���K����(���"��Pd �J�7ݺ�-_:ܧ� ����i��J�����1���QA�)��֛}yuUԼ*�yZ��u����I[D���=d<M`�Qu�c[�w�;85�q�d�{���YH:Y�c)���y�� �m��D�:�aT\��U�vr�%%�ggg�}�l�����L[_�˗��)$EԄn�gI3sUm#�]���,�H�H��,]�Ƣv�d�A���	�b<
5��.����a�v_�kQM���H�ud����,�Ůĥk���B�� cCCN4����CYכ��J�Q���eܨA��K����Z�UZ�|�tqq1�(qGN��c!�p��˾��E産C��* ������C��������<OM�X��rnG�M{��--QMM����

(�!���i����Ec���5z�4J~rʹ�͒:|$�{㓔���N�с#xo\z�!�6�
T��9�5���0��7nެ)�+�N�%o����EJ���XOm����]<��QP.��^9���խe��5ݱ%%r�܊�u�����:�RN��'��2p���+KaBa)�%�\�����p봸�=�B�� �����cW�C�Ҝ�e��l�P��"i�o?�������/I�����,��T�<".�X�p�һp���*U'�Դ�ۉ�B���כ�oF��	%]�H`>~���F��k�ޥK���^�I�̴���Q�%e�uأ�*J],��2�����~u��q�Z�_#��X�Yu�Ȣ@R�}��C�/@�qF�:Ec�k�׈|G=I����G�Xl�y�:2:wZ�Y�*�Cð9�PL�٨g���"��|��B�!�Y1��u2vB����lVgz^�?�'X�9HX,:nϏ�Rvo�tyz9��u:zqF]&w,���|"�uzz:��ӷ;,�3/ف�4
aꋥ��X7���"/��?�`��� �mY��I�F�ʻ�ө�%XHgz1��3C<�z=�������M�/n[#��%�$"n��j�kew^�������X�#��v��8��V��WM�=J:_s���ANV�;��y���>-/.��h�B'�)�� p�t�7գn�UsK����)6LLlv�*��̘M��&;��]��		␨�
�0��aW�.Q�Y�'�6Qc%�L1R�V�ER�6��������CB�d��|с�=C&gg��z�y�������I�A;H�(���r
O�y��	�0l�u�R��:��P+P��_-~�����"ؙ���|�׾mmmZ999Z�f rv��͞�/�a��uV���)@4���.]\@�9����q���]ee7He�3�l��
�uR��������0d�h�����_��}�Ơ~-c�����7n܈����>w�-U/3x��Y��8�h��:.�#~^�ok��ez�L	.��+�7�@��E�ĹI�h+2=���tq�!����+���#��0��]J�?�vHFN�d`ˈ(��T?�4�Ƅ�ֲc�5݈-�d�3�e�"j��J5dv:���$g�"�k���X�p5�,�Z��X�:��!;��͌ҥ9h!x{ZA�C��ސ�ɫ��=hX���%j�	斏Ʈ󉘛���s,َ҉�K㨬�J��F&` �o�s	��Zbe;Y_"d���@�b�Q��0��:Z����An6
2t=O�?JC��I1�Vw+�pJn�l�BMZ���v
�M����$ J7Wo���_���O�>m#�Nʀ��	�M]`M���|��nSDqy����%J5E�2���>��@��Ȣ�=�*�]����_� ��^ֶXq�W$���n��⼁�6���ظE-�Pԉԙ��:`���[YŕBvq����i�<�6:1q�yd��h5�/�Y�<.��Њk6B3n���Y�܌��4 #�:P�hԺ��Mi�L���<�q���[�W��ᦦ��K�e5b;����~�'ʦ
�5�<8���=�AR����P���T��ػ�xzQ�o�֬d��)oɳ1�׸�;�jD��

��أcccr]�0���);˼鸹��� K?E�Lx�9�=��Y�bH��4Bg@�Y}~�����B"��ZO����w�ޤ���j {"k4n]H �Ine�,;	�� B�{ooRm���uxHˍqYwV��`�%3_��гx��FXP?�ۛ�+�%�q����e�Da��z�~t/��L���5�3��>�wtǎLL�[Z7m�LZu�1�k�5,������wd�������)bB���Q�$�~��%����LiN@���^!v@��-��ء�84�;w ��>�F�������Ɣ
:�������/�Ə��r�V2#�H�5H��m������ˋZ��[��x+��g��>e�v$=�8Ib<!�-&&-�:���у^ޖ���G�/Z�63%��R̓�!Z�k��P"{�ñ�4�i�g�S����M5�jt+@�7蜭
9���D�.y���A��ao!�L��|�F.s�D���F�!ȓ�N0VfzL�J:�����B�l`�]w�p�}S�����4�KD�����3ޯ�9F>�A�鐺�ΟgG D������Hۖ��"�qi{����܍�!��jnOv�Yt�?�)w���|"�kvv69le���������q��v ����C ���}�D��0!�v�x"� L�����cb��Y�/�yu�㶈x!>Li�y��%RY�Wx��h�'
�;��Jĥ�
�}���:�Aڣ�`faIҠ�95�2�n�4��ЗH����B��WWø_z����iS4�ĉ�q�r���u�+D��s��c�A����h�KK5<�D�^�=��z�OK�}�UIVbGC�	��r0*3�b�QY�wɲsHX�����TV�Qؕ�Sͣ��U!�]����Ͷ��~?�v���� n����d�P�̑n�g#j����2�d`SI�(��f��o�*�ink�B�r2��܂۶����,&n�M�,��Oǰ���k=���'�gGa蟀�.�vUT��&��X&u��y
<y�%yR��T����VN�}����P�1�1k%�|��46�ST�:V/��ǔA�A$j����2�QZ�&ɁFl��¾f��#�)u��i��K�;�Az6��:�*3�7�<�;�`;3���Y�s���uA(�v	��4�=8�ʾ��>Dn�
j�E)`�|���!Sh8��X����hD���
p�����g6 g�����J�(�k,֑�{�&���e#�HQ���u�� ̻0 �E*1��1��Sh}�wt 5S���q��t��]�J���cSRP��WŸ����	f�:��G�4���_鲐�?j�꓏��L��Gb�uO�\���r�M�)ӄ;D~�	5N��A:�����M��yT��ma�sLj��&�zz���Q��6G� 	4����MN;`"~ZqJ	+<^�r��x�����/���9�pw�qP��{����сO~�AjMMMX�\YSSs���ԗ{����)w*@
Tz��ڰr�R&�K֔�ԑ��fj�DĶ��3J��p��'"��l�q�`�P�|��G�^�H�d�б����ZU{������~&�J��2#���6����S	{'d���?�mi-�#��K���'V�>H23�ۨ����a��l7��DDDh�=����b�Ce1�}��0���^)�G�<fPhݼI�h6rL�Ja��xuW��.��Y"j ��x��2�6J���>)�gQ�V����r�w~�T>צ#����#i�D~���¼���x���w�O�Q�d�Mu{�+���,W�r*H>�� 3��c����
�XY���� �{
X��=�����f`���E� �@�.��$�5�]�TUo����FY��o���Q~�va,��&��<+K5G�rf�vr�{E�� Z���=n-���RSfT��g��!��j�	ʚ~�l
W�a(^ڱ
u١z� ���' �6œgQ���y+`k` ;�F_���񩪪�<��"%kc����Q
�)dط��χ�n�`ع��.��Q�8�8ر�hW���@����
�e_v�
�?�L5�vG��kg��p<b�O�W��5OhSxx�o�F��V�\���<=]Ok�
�k6�S���yFF0%˰Ə��B�^\>dH�=>�j:�q���.�	�̽�>�*�PB��ѫ�L��x��k&�L��O������Φ8�����w�i��<`�8�pSF���/y���Ѩ�J����J:�]<���,���x��×�1n�ŭZ�������A6E<Q2�j��u�O��h��J6�z݋���ݫ(�zO�/�/44�R0�����~=pP�hkadHU�`�Al��Q�*�}  5�+?~\GWm��JFb��BC�Y�.���MX���H9P
����<�XEy7n�hV��Ի��ⅈ���PH����%�S_Q��TJO���u��c�GG���2?(�ߐ�bE��-v�{B/ 2�L��'�]F�`D Ea��2S��pT�Ӕ�����X�3�J�c�~�@�0>E� �P�?<\���������I[J[ZX;��:��DT���C��@@S�%��9�`۲��Rۦ[4V
�	`p�H�VN�<ʘ��{'��c���^�խ���GU_�{::6\��H�L|]4}:������G^�.�8+7��r#�1�݉���ʼ<�D��^^�޻uF�{K�X�	/�L�?�ޏH$�IqE@n�G��!���M��	����&�o�ܼO����u���_�%��q�������$��x�Ow�����W����W�&j�VN@��WX�踞����U�c�8�>0���@�w�ct������7��9�\D��r~o4+$��kAlv�/.D	�E2�hyxx��O-����Yv�T266FZ�1�V@�9�3����&��J��L����IO��5ݔbP����7�����=��8n��-��̓���Pj��l@�Z(��쪁�ch�V������\�h���իW�5Rvya|�8��s�6� �r�Yݒeny�By E��>���V$G�]6�S6]�˽˜ঈp��21}�j�@.�N��Ać����ς���AG�a|�'�ƨ| �>�J~S.)��%��6U��ڿ���OQ�r��Uកg�cD���GI�C8P��P�/Û�/E��s�{�h��c�!v��v�#�N�b�@�no�֜@��9v�9�퓀��� )G5�3�ފ �Da��_���9swf�t�R>�'�)�R*�6���sb����

����&@Q ��8���Vn�X��(K��]@5���mG�g�q���b�{{�o��d��.���uG�ЅW��U��ܞ�,�Lj�B���Z�ῐ�?G'�ھ�\������K�X�k�`���8\%Z;�C�䂚�>�4ee����>�9�X0&$$��=cg����߁�{������î�9��2�{���k� �)W��mu���z)))�0�e0�@�����.��b�e��H��b�d*'Sѣ�O�Ao���	���򳪨���AU�njlA�˛�e\B��_R$0G�k�˱I2�ߡ��+66���VA`y�⎺��.�ꜳ��4�ѥ$t��.n�ߣ�c���:�N�����A���E+� ��S�n�r�b4����K~�3=���/�aFU�ъ��r��-���Ы���n�1�}�|�5���"��Kl>�a#�YhnnyIm |����*t�1E�'�r�x��ȆXH�����B��:thT�sB�w���K�_����
��BB��@���kx�.��R��U�:�mܺ8Љ5d˹���FFF��Þ?��7�.F�����(�FA��ϔS�v��E���U���@G0ԯ� �> ы
��7���6̼��t�ċ��g[��:��k��:Ŷ�J�Y��}���c���'��A��{��7����X	���`0��l�T�%F�P�̼�+1��r��,�T	��-,,�����A�:�42 ��뼎?��9����D��FQnq>�f%���*U�"��|��^��Hq��Rί��ji1�:������L�H�Ofz��<QX��Zzzz�ʅ�y����M���?%��m� ���x46fO�H�\�~ݰ��W/ �(�4Y�4�F?Iыq_����1R���葘E8";c�04�>�+��b��s6ғmvvivew��b�0�ʓw��#���~y	�{86�����u<	>��m����7���}jh�7�l�A�e�V)�#�}�Qt�k�&v�=8�SD04�vw5�.�ܖ�;BJjJo���)'�`����!%�ݽ���=�-��9(���!yd��X�mص#�t&����A�������#�fdϛ�麻���3�S�x�Q���/�H�dmS��wWh+ڦW��]�G6EGI�帖���	啃dr���<2Y����x�	:GV> èV�N��O�H�.3 <ѹ���Tp�'ORΙ72��+sEEE3z��~9�{<��|�$�*UYY��-�t��v�Ζ;��={v�g+qT�L*{�P_��y�a����.�O��	����vS.T��]:�A,�F�NR��qv����xI����r��1���(�u��;�v,�Dw.�����R�b����u����F�G�tK�T�~ѣծ�(��EҖ�����T�/}@Q$��m��eSZ���[� ��3H��H"�4+��.Q��7��
���@����PzKQ���1~aa	ۻ�#���ZN�m5�!��"�G;�
��tZ��_�Գ���w'̍� X/�.N�#�~/a`�N����εs~,�pٍ����j��Cg�讽����\�h�M�A��x'�1\@���	�᪞����Ћ˒���9���&Ƃ~BGP+WFD� :����o� h!R�{�-�#@� F�Q��;�y�P�Z�����D�|�AO�O׊SB��(����h<@}��8nE`li�s~�&3`�_//N+�R��m@���*��U�X�6b%�t:�%5袞��(� �#����r�Z����Zq�P��?�\2}��f9���.��_	���� ըe+����aJ� �|萐xc������G`�T`���0
��T�^�F��������o/�ɀv.G�G�d��?{I�V����ۇ+~��5$�P�<�H^����;v��>`f=��y_y��=B�� `������/z�:���9�Ά]��Մ��Jщ2���gm�	L����pr$����+��%(F�,6����Fm��@�mQ��gՌ�5�/���rFyN$���#@����]j&sg(L��%�&����Ǧ���u�?QeeT��1X���X:�Z�o�������Wj�i�{�Y�~���F[�AZ/����A�:y���C�����Qy�H�cS��y�."��}}}*����$D�������s#<��EZ�����sM�.);��:�D���υ���7I/we��w����G�~�U�c6��~<��z����6��ƛ��C�~Dg���4v�Q[{_�?�o|4�{�y��硭���S=�Mt������M8�Ǎ��$�bZ����Bx]�#��~�ć����D�v;;,�@E�;�x���{"�o3���'c|��i6��&�z��<ʽ���1D|���v�m~}���x��4mL+/�-��k�>f)B�|�� p�E�W�kʼ.?K����$�U-w�����b{'DnNE��Ћ:,�Ѧ��e�Ś҅ {�t�3 *yDA�Mt,/v����Р�ݤ�A�:��������4��*�/��K��%�i�2��өO��a�F�|9���J�Erl:�ҍ��`���:v��A�K?}�">�%����*��!�O1Nk�#�z��{��$3���[�][ڑ�O�A�loLs8�v��L�D0�4$�h@�4��9jO> �]m�����R �#-��E�Ν;MR���ӂ��0�@1����f=�]y4#�X	t�ϳ����������N)(����wov��=qx9�/��z��z��Lt���Pey:�+A1`����s�Nx<Y C�;��[`f�1�z�oo�3���[�n.]�Z�_2O���vb�K
�c���=77��z��_�}�?�؎���������7)������dքH�kld�ϵ�l��!m���Dz
lW7(8�|�1��dV
��޾ͪ{�1*B�288X�UN��X�Ɣ��'�;��Y��_i�ndccs��l1ǽ�o��.O�}������b��6��dv5[f'��2�ij6�2N��=Ϟg_�s���\�	~=�����Uv�ų=QX�@8�䙇r���ɲ�ȹ�?����SH���`fjqqvm�ŋ�5��;�|���v-??�e����� s�˗�X&i"[�]%L�o�Wx�}�I��f�~�z¥/i��p�I���/*xΔs�1�Ӓ�h�lIe4׿�z�-o*�������#���XmC�O�.RU5N���cץ4�Ь��V�Y0�Ž���n�x|zZ��A������w��}���1K���$�o��6E�>��Yv�R=}ݑ&g���q�o���F���4"�Y���N���;�g�����t�u�>ncF�ǲ���Mh_�d���Zi�N�cRJ�6����r~����hwUa�89R3KR�^��5biɣ�9;G��] �@d�B���Ǘ𷈤+<��		��z��uz���Tp@Ȳ��^$�_p�M�q�����+7��k ��q�^DH���"�W�KZ\\<���U}qq��?�h"�b`qM��`zZ��E�_��20�@�ƺ-�/�l&&n,�T�����j�AG~u��器�y*�s���z;]̰�w���XŹ$Ϲ�ꏏ�Ů3�R_K�Ù����O&���rȮF�ib��bbڈd���ߒ�T��0� A����0�q�ܚS4� 4ū�M�:Q~l֭I
� �4ИFdgA��$rt�G�BGC<u.�ᇆ��v¸p����]�9�H�8����X�5��	���8d��[��~�M�W ۀ�����&6�RFaa��/��7��/H��T��񦦦^M�8�M�~Ih�J�d����g�ݡ�Hh���a��{id��~�̅ό=f/��c��u�v��,�2���O㴍αL�%n�E�a�m���H�� ��{�f'����L1��I�s.���|� ��F��}dL���kW�f�ad���Y��q���a�4��=F7�?�d�dD����)A7;vip��1�Gn�DwTB����x
���j��2զ!�tI΍�,��&2�i�,�D���v�Y�ﱕ� �O�m��`[��ۅ�Y��YJ�=�\Br�*0�<p�|������iڶw	��z �%pΗq�mhh�K�K��Y�	@Jj zL�]�t	�a���		��tth1s���!'MLb	�,g�TPp�(7���Q
.B�LG3�u�oJ;g[@��DY��=ʯ��o2��	]n���S}=�j�;��e+%i��Ra�w��v���F����J��C��!���l�!j���:�O,�2�������۷��-����I��)�v�~�)��1��w�d2�����V/���8$Z�̛�2��x��֕I>:|��ev6��M��D���9::�&�c��I[X�8�Q���){��T�cWY�ʮ^b����� �ޕ����I1M����o�U%���y{��� �y�<~�Kέ[~���ӷ����@2�yp����7LT.����_D*�D��g.���~�g����1S<���)[���0}�����e�m�[���P��8~�̀.I����#22VT���	���132�6Gv,M}����*�㘽~�}VZ:]�+CEL0�H�qƽ��T�S�y�i!��|Ȥ��*�v�â~�d�ê�<{�ۣ�v����{�fY�@�eѭ�[d�u�s�1�,�\���ڎR�[����|��K~��xmmm����ׯ�2*�	����L���{	�a��5i�1����i���*��m��~�E��o���?iz�m�}(Z�]���CZ*#]e/���I��G2� v�DS^I�2�{�n��ӧ�B@�R�����9u
�=�Y�1ʦ�^��IH��D������Z����x�@�]iLѥZ�ʅ(	��o�w����4���^�{�QUS�>~�G�e0�V��5U,���6�i@��[�ݧvĢ�s��UP@���.h���տ��p+��!��	w�ڵ��a�%�ג@�#�d�t����2��2}?~���ƀ���`~Y�i-�)�7@�&��Wo�VE�[��J��6t@�����yрf��e~7x��5<M<��=h�{��ly+���t��� =��mbB��6��(��~&�g��
�.�=>��m��}l�s�Ƥem׿��"��pJ>ML�dp������Qq�%�����@��l�/�۰xy�v*��ZXh@!�w:;�����8����1����f�{IK�hJ��˄����z���'A�׼���OHH~�ܪ�ȷ��e�G^�d0n�Fd��.��7��l��عs I~1���ð
��{Eh�@F UW�Ux��4NG��A(��[M�X�Ƀ̄����Y^��-�J%A�U�jy��t���x�c��`��,��bbaa Ȥ-����|�P>Y�r�wö-ws �r1��3��z3��у&%�����������k8)H��Ѯ�q]�K�0�ͳ�9@�x����`��V�@����QU]@P0��+ `!���}���?��4Uo?P5���b��Y`�ɘЯ��H⹊�\�^�*��x.!!a�J���&���
�A����EkUqpȖ[�1���/z�1�"�b��?����a� �����{6��*�����}��s�U�h(��0F�p�V�\u{u��o���ÿ]�_�����?M����2,M�ѵ_�_Q��jaٜ����(0�9>�q~��zLI��_1L`DoJV�G*�T5��%��F(�'Ҝ�&���Ǯ闸�g�&��'�I"���_��6t�c��q��*?Y��+�Y{ěVYhY��q�s�˰��ΝsY�퍸��6�[o%J�HJ>oLՃt�
�G$�l��3��/$B��%���dΓ315�ĸ�7<�t��Oi1X��Y>$���V4���2�)�UG��I��ЍQO^�� AW~��.+�e��a�n@���/.��B�`�QWW����؀fF�Rwlp�x���j���d�
Y���,�b���l�C��끙'�g�<���3O������qtI��6+���~�p�Sa���{�8l��r���u2gv�����������-Tɚ�*�7ک8� �}�Qf<vd=H�4���T�#7�#� �+]�a��v�ݻwG��d؛���$ &VP"���4��*M�R�����87	_��X'Z�}�į�l���1�O��t,@��x��n�s�Nѹ@��z�h���>��$R��jH�;}�=�Nd<dy&dŉN�l�]�	�hT�.:G��a�Kc���a�g���Z��M��g�StS��Q=�w��irLW@@��M�������D3Z!;�J�Yy�U+AV���I��s������g��	��m*�A�]�e�s���X������Ů�����֛�S�>���;�ž�J�TDYCZP�d	�-�ز�Ѧ��&Y����-�#�R�PG�Ph!��?���������u�y���y��k��~fZ���<�3�kr���T��l;��o��ߏ��Ղ�������0�枚˙F�O_�U� x�V��RV�	.6/9�	>�G�IJZ�@��xɋ��o�u��3��sѬf�?a�����^!�����	׃���ij���U�x�C���9oE?y��*�0l�t��/7���Q`ᓮ{>��d}Xe^DI�a3$���dZ~�:FY�#�W�/���나P�[����4��#_r��N��S[���%-��[��%�o=�{��?m��9���ϐ$Y�G���{���;�������7�+N慞)�����)����c���p����D���GC+׮�{�ҵk0��6E+�b.b��Cs5/~$��[,d�C/v������k��}W�k����ۖ�R�:��s�������*z�}�^B�IFY(�F]?�n�rt����O.���0[�ߦJ���mlh�˺<==<W���(�꡸@�U�菋7_b~"��6�RG������$\��+��~Z�IT���I�T|����<>O$w23�s�, H0l�Ѩn�A�Ӥ�sqr�}41�:X�+6��G̷��޵.�"u���6M�z�bbu�E�n���ih,���>!���ϗ\v�065�-������}�����5;"�Xk�jr�__LMҜ.R�r�|�s#�H�<s����n[�+8�� �yp%�p��Ƒ+�J��K�#�:r��������lB�˺�;s?8����	��<��҃׭(��~,ή05���D�.�s�� 8�X�_��Xtf+>���ߴ��G�
����_��;�z��Y��	�(�G��T���F-����)��]�&:r�����p��j����@�����2w�-#��ѭ���.���5###f�����k>�_!W��K-U;��3`�~��#�_��|Ω�':8,C�

6@���E��R>�[��f�9V��Q?��adj��7L�[[gc�r��f�_�2���O��5����P�����毚���/�6��u���=���Ϫ���FjEDD�����0���NP[��� ���r�y�,�����.����b4\�|�l�3���;fo������4��l�k�wo�<GG�)��l$<���?��9�
y��@IR�������߇r'�����gՍ�����\Z�J�Pk���0��nnYR	��$6AN���~�Q�
����u;���]01Ȕ�n��D�7�WR��&=R���m����|�Eꍐ��DB
�0A1���w%�
�*{���H'B<�=<��㋄��Y� �w�}�$����;�\
Cd�Y�[X�||.4�I��d;��m�����r��Z�	)�!�eʆ �x�G��Ā�Ʋ�FT?� I��ם���1�շdZd�<8���م��ѐ���	�˚;�y�����7A��f'������/p����>����ꁘ�����J���LW8/��EQ� ���o߾v���D��4Z(���V�`�R"I�~��_�1�����Ɯ}率K��v��+�ظq��o�}؆UH�M�ɑ�\���Sʁ���:�N��C��g�8�[b�ns�˚4�`�˗{ �H�ϒ� 'w�8�|sG�]>>�$%�֯$�g���i@�?�c���Q�Q�D�qX\�����m���@3�ED�	'l�ܖiII���� 'e#G��ڙ�����GMì�~�{]�,���+���L������\}�w;�����x8N�%�dU��]���Z��3<�			Y҉A��,c���J�>;�{�)|��A«�p��R���o�[�'n�raQ�8'��K����J���V�wy�'�َ�_�*4ݻ��fZ[W�w��(�~�r�����j�A8 �8��V�	~l/<�ui���f�����/����˖�kη��x���gq��#���TY<��b�������\ s`Z����Q��`do��9�/�A�Wo]i��S��*t���*�.����gϟ�|mN �8�����1��������c��LDm���U�.:�D+�����uu��6O�)a�#����a�X��� Rx"T�
y��	ϴ�XS���6���Rk�s�yc9hm=:*i�
!�@xq�������|;����g|�㟜����#7�����Aj!��D��l���9���{���4��:��,8�1�	���zg�;Qc�?67nm�ȫ,��_��U��c�`z�azix�+/�	�t��! Bۥ��J�*�~�T0n��u�~-�ɐ����J�b�iچ@�m�sihmy�|6o���u���E���ʩ%��+�n�1[J|�
�u��*\v���_fuD�8�^��K�46�cW��:�2w�#�����;@k���"��>���;w�Z��ܧ%�B2>��7��M�W�޹��wA�elf�}���\�!�u���#vg7� >ڛ�L˵�$'!ʹU�b�*�N��� ��e�#o]�����+�:�<��'�<��8�v�|�~�j
z�%��� }��/���]����U�Dc}���oQ3���>������.��z���U]g��Y|��E[�e*H��>�Ƈ�ԑ�]�l�Q�>8	:s�|�O��I����~�q�����n򠾎�a�+XT~��'kAjj�*S�л�[��7�u.��J�һ0Ѯ0���<2�⣼�$ �h�����4�Ʋ��<R���1`㕕�w��%OX���������?K������ �/���k��z}ĭ�l��qV���;�*�Sς�j��t"Z�ќӾ�m��� �������#���J.8�������\��odt9��c˖-w��[�����!77ܠ�c&�UC^Y���葿��^齺�DR �~��-����6���L�V�A}�ͭ��*�>|�xhr�ם�,rwVx8�IQGWy������]�bϧ��q*F����QL������CA�v*Y�9�;w�v~~�jy;XS�������	��1V!�;�F����V��^\*��@Bn,��o�"�uiH��\V6��ikk�U����1ɹ�=�P�U���ǻƳ�4f,�	(���3[ݓ:�s��i��	| Jc��ywn߮V�[�:��K��O��|�X�h�Ft?Y���Ĥ4N���y�֌�#�0�S��?
0quu}~��V���Դ�H�W��W�%j"���I���o���|>�tr$;���f;�4���B�DUU�+[�$nܿ�8�H�:��pb<��H	�qrUD2�����O/�[�f)mؐ���*A�;7on��/�����9��L�������M뙳�{+d}����ǊO���+��L�򙚘�R� d������/G��a�7����(������6_Ȇ%��ԜZ2>%��r��A�����2Ѫ<^����l��n<�<���������{V�6�|���Z��Q�%������j���e%m?�;'g�}]�}�ߚ��ys)(%=7��!8���s�'h�N������l�`6�:�q/�էDd?��?Tv���ݻ�G� �W���fw�3�t2�����d}���Kw��	�?̴���?�����k���oK|�!�^�v--.Nt@�VQ�e�Ye�%"����L.,4el��d�fC.���Чh�����L�nMN��Ȫy���߿L�ulP�o�����K����3��O^M��O}�o�2��K����̋�	�&D���kK�o�4���eN��
[p-���M���A�� `���ANsi�r�<l��4ѽ��*�{����k�e�'����ۮ��ד�w�����|}Uל\\�$�qpH��'����/�w�����hbgle������'q� j�AII�w/j�� ���e`�u���6����SQQq'=R�b����7SQ�����	�5��f��~�u�4p]�9)��ش헥��ʖ��~����YS��6�7�����ϱ��2��w�j���in�HJ������`H�����$<��(���|w�K�'��_`���kͥ�0C/�x����C-�d���b���q`sCÍK��ܼ��ug����������g�i �1�!���H�Qx<���9�!c�;������`]"%׳��/^��d�	����[=����/5��B�����o����;�����2g�rI����><�����g�r�����e�VJ-�o����@��Q��c7|8(U�E�>��K��8�X[gǫ������塀�����f��m�%�ȃ��Pu5*��o�}�L`,��o=LJZ��ڊF�|�����I�5�#�!We�RZ?�>M�tUwk��Ϡ-eH�1����+R� ȃ7�⮂z��h�"A_�pA{��pE�ɹP5Øne��[r�j�����'�օ��)g�E��p���[���K6�[�]Zj0h+��u�2D���K��\��耬R�?��N.A�\ED����bbc�8�L��Ib�ǿbժZU�54�?���=�,��$�q�W��	r@�m�)ɋQQ�ǎ1ÓkTY�;�&�����}��SU֢e����0��<�4�z�W��ADt��O�̿.���,����/g>u�.�q��dWГa��OODh+�=1�"�_2���ᑃW�q�瀢� ��[���`�#4b�!i��xzz�v==�ւE�?� ϓ4�9wm���f\�;%�&O1��E�D�܌��GYoW�9 +Y��Ջ� D�Ǝ��*�����ھ8u�FU�B��̭���Ϟ=362JvnJ5s,��$���de�G��R� /Z���m�D^m����-s�	<]�k$����5ı����i��F.M߰u�E�3fy驩�)))xBə�d��9h�!��������̢��b�u,�d*b����f�҅����Up��tnTlr� ,�ML�b���ۼT��#�<n
�x~]�e�N�5k���Ӌ ��7R��b��V�~�������"b�5�IL_g'']���vo�~u��z2�H$������TTT<�L����m�S2������7y��<6+D�]��@�3ٶ�$�q7O�)��<��u��q�j�+�s�?ʆ�Ĩ����w"����EڒP�P��ލ��X|o���9E��L�H��@��,�K|���K�w��?m!߱..B�R �Eݭׯ_��z�~�
�r��I�xR������p�ӈ<E_����08�k<u��K���F��r���t9IP�=Eu���7X 
�Cʻ�?�̑�������y�Gw�cy�g������[UK'N����Ͷ	�(`Ïϟ��i1-���ҷ(t313�ο��6�Fs�q�v�2�8L�V9�+Ʌ����_�ƁO=y�y��{ZW�^%ώ���9�	a�᲻{1y zVƖ�;�h���׫W�RS��V�r8��ڮ~����������ny�֙IK�X>��6����?";v�(�4� ��d)%ʭ�8X!��̥�B��?oߚc%K0-,�R�d�
��ۜh�]^�5`��x6��$��]w��E���RJ᧊t}�y��R���u)�ғφ���������D��b�Tb}h�C���`�-���xYڠ@��Mg�ˑTކw�&�3���vH���k�e �E��;|�i@��׀)"��$��ϫ���\�� �m��'d�xpZ!rsVi����]�G�W�̲e�/�Ф�����׭���a��q�	d�O�C2K�B�°BC�<w�&a34Vœ��"&�0�Z���\,� �=�g_��f>�,�p�Y�PɮY��n�FFgH*���X�\��o���E���G�JnV6���d��ITrK~6GFFa�}�r�����!���\Z9����,,,o�d���FC`VW�\!O�u�Z"�?�\<�$%�;������H;��l"������?u�aA��b�/^p�G�A�� M7�ڌƂ40�/�W�Us
�W���<�=u{���OXy&�3eٵ5���͂(���4Enɴi�2�	��Z�����==N�t���g��Z�ǅi�I���rk F
���;�
%�>-�]Y����`�J~a�E/AY��Qܘ'g��Bۜ��X�����5�,<-Ԥ��A�T����HE�����5Y딕oi+̀���� ��I5]���+B�iw��'�1�=�.Ϻ&���hXg���g�n���y,��7�I������2�U BCZ�����nU�#�R�mʘ�MA�kq��Q>�[�K��a�S!.��򗭯mij*�b��sf�ׯoWVj��� �|������F��qk�	PGk�EN�����\�
�@s HO��L���hl������M�]k��������P,�(e�2>��C�28]�@���b��2��7�<0���rN�<���Y���>>>�(��
�!G��C<�Seպ408���g���e$��gWF�~[��P��y��ё�+��Ő��{���(=9�B�/}�a�����Ԕ!���D؀�z�,�nޢ�����o�ۏ[y���@��٦t6�����
���Bƍ8�бS�[2\_��[_�!: I��c˳n��'Z�� �1��QrO ��6,��o[��,��]��ѣ6"�����W@`�4Uǣᐴ7��W���pOv?>��Ԋ���KT�,F��E1�j(x�U<Z�Қ�|�K��v]L�z���O1�*o�8}����]o�n�0V"�'��B��W$�x� ���
[DeC��k`K+�s6F���~h�;���0bH��CLv�l�ڟA~�@n���C���zc�N�B���ooAp����ת�� �C��J\�0;���W�1�n=�=��b/<� ,fd�|���}-f�h�,���QB*oE�������lr�^p��9��ɉ��!!�DY�Ǐtď�b�t+��j�X�=� < o��X\y3�������*Տ̧�s�6 	*d��m���ԃÎ�ơ��^��Z��E���ڀ�{���OD�V>��}�ˀW>�����9ŏ���;��-����?0�pݬ=�������ON���̿}�Ύ�ܝZXh21`]|�Ӧ��w��'�����zEE�c,Ny�`�ʌ�D�km>����͛7�F�������<�ܲ A�m���[�GL��:�!'\Pa��x��$9rY��Ǐ�̥�R�]�����H���x~8�8�����	&�&��ǿ�9m�nĕk�/+�q*^W���X���?�f�Q���#,$�G[����.����ߗ���x��� �l�:M�<���6$M=!"*�
|�?G2,�.L��	~�W\��#��Sz�L~]#Q12:z1&D�f�+c����m����ݖ��P�N����e��A�x��9r�ѣGQ����7�����!��� ��'!w����|�E�����),�OXke�eKy��z&�ޯ����)a����9��^c���>^j�03�~�����Y�Z�u�l�w.ã�<�ٌؙ>��X�lYuA\�'�r�.#��$�5���������̡Y\�����ލ�g ���� /�2utrbN���2��,�
��y��
�qtt�Cv�����'zS����p�O�h=]a�!��o]'����:_C�4�P�R�v@&݀VM���۠ڐ]ɛ���ޝC���e,�N��N.9��1>����x�(��9Q.�k�B?�m窔�#�dN�W����Ct̗޺m�ggƸ�I҃�W��cR]����Y����|�6�c*��M.8._W������%KT�75>	
�?�iR��l�uy��j_㇂��
Gww���V��_�Sg�'��&����0Ǆ���fkx��y�t�O�V���{��c��_�{�Gz'>�hzz��l��,m4}�@�S:�Is���~�]q�?/�A�E�)���J��}�O�##��Iˈ��ѹ�lm�b�~�C��{_��J|���9c+Z��%�i��2�{ڃ������X����`B��TI�DV�5�u��IB�E�����x�~~�J(2���6Ѥ9a�]ݱ47]��)\��Pk #` [�[��m��X�sj�g7���&����/�����/�Z+Y|���<e������S�X�Z���H�W�<��D,}�?]��BԘM���!�ZQ���|+�b���j?�d������H�Bk9-?'�9�������A�)�i;�V9�4�g��QOu��Dk`���?�S���a��^�|)(.~; EٛNkN�`�_���A�Xק��Goc�CL����u���sm�������Z\�e�ݿ����`���X�ï;;�s�lx
N�yf���_e���Oה֯���-�
d�������� �0L"2����ã�Ѷ�X�뻡`%l�����p���*,���ӏS>@�ߢ@� eQw���i%��,�2�a���Ԛ�~���q�w�K�v``�8�A�W��SwRۑ���<��to�av}J؛��2���S�/�!�v#􌤙,�o����1�TG�J���[s��4r$�N���_�C�b�)fMg���^)P��H�'��3gμ�Kh�8ƨ2B�a"�\��q�RҤEq9 N��Thm��e!�|����Z��^S/�lw�f�9ƃ"*�`��ttt�p�\bx!۠�*��g���?c�|MP/|��G$���g#ӵ
�w�Oj�k��⍱����L��ze<���\Ƭ�E�k�A�arH���;�0�i����Jh�qQU3�=˨\8�i�$}���Y&��^"����$o�����=�j%�qH1�`o5��|�k��^�>uU�̯*e��R��1�VvEU뤞cL"e�{%�&�~�)�C8>{�g`&l ���5I�i�Dԙ��?2�'{d�w�~�p��b�rFk�l�	Z��xç������a<U(n*�o$M�+>��1�Y��E��
�������+��d2��`sxC�Ŗ�xC䎔K�Ҹ����5�.�C�N�! ̍Т�B�c�A�l$,�,��$�kAK,�Ԉ:_h�y�I	�ʒ]s�@�rӜ����+�LYմ�v�D�W7�� -U^���K���"8���tV��"N���rD����_�`w0݄�V:�o������2��;	j�`+�ǵ�+8����c�/YZ���rB��Z�K�~���lD\kK?6jR��k����+=f-�6���JX
4p�?~�������6t}7�\&��� ��y��t���U�u�����? ���*���c�W��v�^R����*��=���c�ب{��;����b.ChNl-��ݔ�j��f�y&�YTJ<�
v��݁�{��3*� ��'s/���$_Vq����O�J(��X�OIS�8�����L�̌ցt��fc�IA�"m:^6�(�ƎrbA,̚�č�uww���`�噱;v<����bߵ�)uԌu�ηč��;�_he8�"δ|f�ɋ�f����R����O,��b��F�ϬQ���O�$ު�`����w+�SZi�&("�t�g����GP6j���q�ꆏ����U�!0J��Э�:� F2�Ak@XPPwz˷��al1�3�d����{U����*�|�yl�ڋ'�}��,��̽�V�iӇ���<����P�+!� *>!!aŵZ��죔C֫��"�g���se}�,y`2ҵ�����♈繬��ò߉|�z�I[�*e0��!�ρl�����#�x��9���Ǝ��Z���%�i0i| ڕ���gdx9I��Z	E~��Z43�n%k��M��+ ^��9i�)��0���/��7Nb��0gAmijk�~�05xh�J����ʊ u�O �H�1�	=`�~��4W�:� ��Ev%{�7��f�q]k*�m@` �<�:ᒃ<d�Y�$Bn������y��'�����-^�v��j����iXrk��e��=��
�k_kA�� �mDg���Ֆ���T���Q���szPU�P̫nn7�����j�� $:se�LO,|۫�p�4Y9J���e�5�ˮ�=�t��qF�LWc=Ǿ�Rt��k�[::��	�!���	�2�s�f���zHVn�Q ؙ�r��(�<�c��=���,��		��A�,Y��bG��=?<��b=g�;�"��I+��vދg&2Ņ��LZ�>��:h���R�T�5��ʎ����9�Zq�:{oFL���Q��kK����G|[U��3����'�V�E��^o��]�yA����%��ep���~���5�"w&�xn��BEM�*++��*���++�t���>���V
[�����hG}N� �Vj�����s��s��/�z��j�ÇeQ~z3�MßBBBH�Q�aXB�(D�|���O��fDb����[?O��f�w�t)0�mϋ�V�ӊ�kxѓ���H�jg���2_H�!,"��c�e�Z[ooE�v^_�g�Y�T3�2}�:|7v��3��@^�����=�v��L~Fp�nan;��CCC�߸���p�m�ņ�Xu�׊	5y�dZ\�Q�ˀz�>4r'Y� w�0���3)���G�	�/�w���[����@��C�5,��Y����&@��z *˴�/~��y׌�v�2�:�`%4=
!�n����*B1�g�e�/Tg��B������Z�`/mpk����[�2��G�P��B �~�h~x���S$W���p��niQrĕ�����x��`;v�	�����C�3 �;���.�"���'ѠNV1�&l˱����{��9�^gpd��n�
x�	v�gcg���};��w��ࣤr�\��<U [��qq��a,�����a5u�ŦB���8����f�6�L��s���
��7��2��71�N;ԝ�?bk�Hql���X����ʈ�6��z��1'D���;�V[ j�A���ͳ�|{��`t,����l��c��y�dD!�Hp�������f�n�� �/ 
����b�NZ�n3�l�Ś���euQ�e�h��(a�� E�Xy��5̀}���P���B��c{�����'�	`�T�8$�?�c#�S\a`��5vAA�@��Ǿm��a&��1�م�J0C��K�9ۻX�c��H�ӟF���&B1
���n�ʳ��c���J'��B����GRٺhZ��:~��)�
�]�v�3R�ՙ`u�m3V�x����H9,�k��5Z�FZ,�a5���dBA6g�.��
�#Y�[�}^�q��:���r��)'!��������������h,܊�Ϝp����#Ǿ6
����� �+��mutt�F��8���
��3N�f��Ԩe�>���J6Lr�s_���M�'�Q�2W�73��P.NNl�����V���?'��m�"T^^����P�XvycE�ɪ����Su�Ũt�D�`�&^��+�Z�m�\FPo�&qU��xFб�_=ܟ6�`T����us�l��6Fm����𺀾xx÷]ha��?ݓ�̫�n���׶��`����Y�8�aI����ྰ���4[q��W���mٙ!O	[��N�FZ�v�e81�����Y��1ܻ�^��r�����S��p)l�3+���dyE�+p����w%���U��e

��p��S��l�f>l��	+�Y��R�"��:!�F�)�k���:)Ǳ���������m�j�m�J��l&"�>M��}�7


�9$H�:�P�0Ya�S�	mq�E�v&� ���h­�z�X�j�n$�H�	 v2V�D"Jjj{��5�gī���Q[��K��	�w�bo�>Lb�����`���-+�$��ͪ��zS�-�?��FivNN+๊�؁�FӚ[�v�;+ 0<8�B��=aIm��_�JN;����:��h��Q�'#D��ɐ��&&O��hT����tEEE^P$JX 9\dL;M�Kd���K���1pF+r[�#���-w�x��M<S@��j���Ә!}U@7�:8)��4�b7�(����h-� >�	����qk�oΰ;xP҇Mq`d�K�]�^y��x�����HL8�Cv]	Ђ�i�s+�A�A��@�1�n�2�<�(�ܵ�e)j�ۇZ#G�r�D�r��-"���s��It��֩�
3X�g�uWyn$	��-t�f���>�$�\8c��~�������]Re>��~+))	{�!��߀Φ#*cl��=}���6WVc�� ��zʎ��DO
;�Y�oӶ����^�0�3����\�|�5�_	5P8������#�z.��g�C*~��Q�?�O���z�G6>�j�bK����B;ʽ��j@��A���:���wz�Z�0x�౮CT�vtt�ąr�؛\�) o�'l��
���[ɗ�}��ϨU�iǣ@�{	`�
Vl�	��AV-�qr3vnę3yY��O�3�-H����w�X vU=��j�	Uە�6	��D�$N�H�՗��9�a�i\� H. �,  �)��F3�s���&̟a��֬��7ia׆-��w� ���ᪧ-v�255��&���1:�G�V�����ؘn0�������(�t�]`H���y�&Ҭ�E_�~�Ƃ��틲��oJ� �[R�b�GY�����ts�����oǦ�e"s�>+�9Q�f����23�!�J;BJL	�i��s�:��O�GV3��2��`$�r���*�p+�T�еȥB�KԚ��d����x�!�`j������!�1�
�>0,/�1��896ޫ)~�X�ts��������lق��Ţ�$S�2��=fv�����h�M� ��p��1�M=�4Y	�WX����㕭h����#��:2:px�k����o< �E�&ȭ��dLz50��72*D�W�+�H'z7�O��E!�׮i),�b���|ћ��%Nd�(�X�N;	~�_����뜕����1p���se������ p��h�އ�v����|�+\zޖ�oW<�^-��D���M�H[?��f�j0�zS�~��j�� rlu)��%,B��='����ַA���3�B�Ug����?��9����g����I4'�+	�ɣG�<����y����K�������1֘xm�w��_p��ޓ�w��h� � M�¾�I k��l�VN��� ;����	���y�=���f��MMN�+H(�ps��ϟ�c��u���h�1�1$�"���Ò�3S�C��<�b���������ua�	�cJ���t���ߐ��ERHHֻ����̹}�������3G�?oq�qf��@�1H����q}�z·�)�f�8�^i/��`:6��U���-5�6��&�/���X8ۓ6���X�ct�f1�-ja��%%�w�=ִH*����uv6B4���L:d`F=}cA��	~���$����u;��,Ì��pw◥����5�m�g���`R��NΜ�����dQ��(al�c�]��y��ͫ��g8
���� mX3~=}�t��A/y9�HU���»Ӎ�b�Ep' rs-,�����Ƈ�Z[����%��vN��~����R�2������T⹨�	�����ۃ����z�!G٨��:|��,���0e�?�5E��΀�0��\�����y��11���1�g6bbD��-����d���0B�9h�o=�D�fv�Z���X�{��(��\kjs�����䛃PY��.����w�4���=���Z������([:�}<6��>������[�Ӵ��E���b�J��oP��$��Bü�R&�+^�޽{�>}��~��݃f���۞Ţ��1_��El�η3�%�}��+��"���tɕB"�{��tV�<g�s�;� �N��7��k�}�.읁�M1�ZI�<�������V�'��1�71�#� ay�Ϫ�132��`s���^/[Z JP� �D��s��@L��K��},�o���g39���j'���q!!�3�A`pաء��u�ò�,I�!�T^\���I�Ý!���o�r��X}�֍3Ww���(�D7s"��F�����[���#���ۀ��8�h�J�G��UL�HtF:�4"D�	�� ,�e�����\YlɊ��go�6���q�ĈpZ�s0TAHÆέr�56�	Wc�p�3�Ȼ<
�kc��ao)�O>l��,��g��e[��A�l����ӊg�}	�]P�<�Ӳ� �:��e���$�6�sr����IWά�9V��<0����z���åd�}`��އ'�f⪦-�����F��J�Uf-f;;�AV��|�u�aXƙ{�S�Y����z��f��"�X�Ǽ�`V�� ��:��^��b�!���b�i6�����cSv�#B�p�<8�mH��i�賰��5׌�-Lk�J���^����Q�9����ʊ�l�Ӂv�}�V�y���$'� �ʏ��(.l�bx&Y�����Ǻ°�i�5G ���ʿ��B����`_Zƽ��2��_�V��T��hF��ꂚG��t��ޕĮd`�ب�\:�>�xrrrү/��M�t��M��z�?o�!�f]U�Ob���0��߅A�������bj�w_�r���Ǚ�̫�@� �֊��K�ut�O
X�&�m�' q�&E��ܩ��P���^s�!+{�p�ģ8X�̜���6�3����2���@'d�>�#�9՚J���{�d[�]����gk8'�1@H�!<�Z,�#�Q �i�q�/z�����ζ�h��|�x��V)\w�a�2�y�=���X��b��ꆆ�$4ҍaTJ `s�?��<�
�{1�����G����x��C��{���y̆���/px��Uk����ث��z�77fgY9Դ{��E+�[a_��(��khL>��fu�V���_�o�0�������C?��G��4J���(M�⺂�Ʒ�Ko�{��gZ����"�:ܲ�Y]�Rg/��bUY��\�Y�?�T�_�����iuLN�Ǐ� W�ip��y�)i��gx������`؛<��}M�**BxԨ��F��o�85�5�N[[��O4��*�2�C���L%�ōWg����11>��ގG����/��~��^4&�RP�9~5"�Z��&��e�Eك'�^��m� �>P��_���9rD�>�м��7/djOˁʹ�NK��W��*}�n}
V߽��׎��S㣅�z�,��h�8fH��>bӠ?�S�O�&`��zj������\o����nę3g�G��׷�RjU���l?��.-��qr/���(� G
S�_X���\�Htl
X�Ǻ����"�=w����0�;{J�n
j���x�\���
�2@Ew��ġ�/.��X�.݋0�kL����e��7o�#��<؛[��M���N��?�ǫ��yvt\���3��|�"�8��L�|��t�@xż�)�޺'s�]]��<�
;����� �h�%��rMUa��+��+���=٭ ɦ��c�;::�F�M�]���?i���V>����B���t��	���vUҏS^X�������� z����Z��[����x<�Ss�t¿� ��>p�Õ�����q?d��S���u�+�؁��+l�'���j�s�ʖ���=��I7�
��z����{R��"���>�!2Pd���HYq�⏄c�N��Q�kş�RqD<��ӧ'�Tk�4���.EW�sZ���-�>�a�� �p@"�<�# ސ���޺���,Z[qG�*�/��O�/`��?x��5��i�c/Nn-�w�0b���~��@��!���q����3 �x�u׮]A=[]�.t$�=�3hb	fb���<,��v���|@1:*��+[�x�>�l�6�
��w���^��Gz�m}
�*��@�)�t;j��w���G�Ѩ�@w��$�$��ȥ#�������@E"~v�h��=�z|�+ׯQ�Sʒ����!��ޛ����Ii�b�yĞ���,���X�k����!W������N�gO��ѽ4B�6f��d�$SO�+T*���;֩=E��[vD���Z���L�Q"�!_�x�/�Y�w���Ɨ�w�i�Q���W�~�J��C19���Q^��ٱ&͉&e���@��o�!��ʔ��e��
"�YH;��H����@K�6�\�|Y~������	։��⢢�z��ކ=�������̟,�m_�]�7'E�;�R�>�*�/�Rw(k�x��߿�G�UVV�����
o�7-=[�0����py���c��F�>H��X���hZ���ʿC��'��MX_P�R����z25�g���J��"7,9@��G��AQ[[�����x�l�hS��]��J��o�@��!P�79Ih8u�'*8�CN�ih���)����p��C��4�v&Sl���=��8nȼZ���R��7&ዀ�!��=>�)�L��J�R�y~�O�T�o��t�џ�H�xI��y9���x/�`�V��3�!M���gv<��N��U�����
��m�U!�:����j�>W��9gqK��ʹ>��˅����q������\�m�ǰ������v�������C��)��+1�$�cw/�;9k��� ��~�냶�Gھ��{3P����)�oT7�U������Z���6h<�i��%���d��ǚ~�G8���+p
^�.��3�ߪ�b�������7�zh�=\�c��={�<P=Y~��Y��q�6��2R)���D��8��Zc��>^��#bu��}���fY�C^�����{q0BK���'�C���$��}xp]zW�.NN'oo�}�ҍw���P�����mjo�������6�����/�Ic3��;wd2��3=��L.���CP�W��;&�|��X�$Q�����w�Ը��k�b�v�̡�CN�3�Ni&��
�,D%އ�L��w%)�
e���S�^<�BQM-��I���ķ�뮿z�:ܽ|���e�d��Vel��FAN�5x3GS��@�����;$�zA:}���O֓��8�*�?E�ˍ�u����7�����!������� �޾�q�\#��d�����o�I�{^�x��rM���P/e�T�,jyb}Zc�!$��9���I�l��0ܼ{�[�������h9�ʁ��G!M��V�K#��ŉ�H:'G Y����6P�zB,�|%.Ж�\�?4�J�� Y���|p���1cu���ʢ�ᇅkך=��`@��g�AOOC�_5�rr6 ��({��m���)4o�l9m1�V,I8:j����E].��6�� ���C �A 8��P����e��W^�QS���L[|�~��=E��H	��φ1u�o�2W��C���x��x���X���D�� ��� `� �@�z�Kk��d�.2QQq
�Trko�w����_���(�V�D���~�F`��͇2�T�G�ȶ���}��.��̒��6M��O��=�Ѵ���e�%v�\���4����*��M�\6x��C���ܬ.�!��{f���oޘ%������XZ�G��L�G�b��q)<�+�NMM�US�k�{�Ň� T�-�<�GZMfϺ�p�OYA�~vͱ��o��Pm~}���{�+�z*,�/����{�/��9����\sBΝ���dne���Շ m��{-7wh���,*���܍����s���ۼ�4��Ws���o{|d����c�N=R�f˅#�\��jdd4���oP��[E����o�(�K�Y>�<��ĥWw�a�2��|��d=�իW�=���M �k߆��Vbk�E����/�o`9w'E���ΫL��[S!��n�0c�F�
M��@Ugx��v�k�?C�#�t4/��\�
$-�1��l�R��6�o��b)ؽ�V�#���ۚm������
b>�}��<
7��TZ��ԇ%r||�cbb���<y\-611��M}pjN�<���(w�s�$�P?�ɛ�*
�E��Z:�a�O_�r�l�:v<JK�1�`��
lnmM{�rϋ�ϫ���e�c�z�݋NQ��o�1�؛���e��w�#�;8:�hN}�<���9�8ٗ���<��o
2�	�|�W���D��Հ6���@ �c�����哓�.������D��gVev�(��{�\|V[���RS��-��e�үk;ӛb���&�/7g�`?0�� ��'��6aϽ��։�������Z˗/OŕS�򋻤|F�MFFF�mm7���3��3���Ibu�
�ۯ ��.f��͹��#Oߺ�����,]I[��`��5��n� ������].>y�~��T枟F⇂tJ|�6��P��.��+�k����k�^9r���{i]���~�"���\Ǔ���1�>����p��E[�43���Hi|�*����A�azS�LV�%W#�+ tJJ��_zS�'D�܊�E���r��bq�;w��ǽ߾}����R?P>>�1���a�.m���x"+3h�~�n!����ڵ���^�&��� ;��/�~�d�~x�(l"u�l���#���|�R�klhx|K����C?E��B�w��7e�����ޠc��M�4j:�i� ��� ��$5?   !���нշ��~�㛚0���P��~|>"��WH ����=����u�m_�`d������X�v�<W��-�~��/�&Bb;��Fl�g�w/�;�P����~�
���δ�����ڌ�/ޙ��?8���=�M޷�/)2KypS?��s�m	.��������U��oѪ-[��V���pD�}i�1PO½�U�S,���s��X�m�֏�@/�c���K1����F��y���Jv�x�[�-Փ��ӬT�7�����v��I�}l3��G#QV���}8Nh[�9D<���((h�(�L�-֪���oT�WO���_}�o�H� wT$Q���~~�j���"~u�qm�t�~�:�F�������;��6<�����lx�U��tYi_�@l��=�reAs j*��.ޟh^�{'��'��7���q��)[�bU	��(wۗ�5�4�nQ�8qJG��W�үg��A%&��+�������C�N|�+0�Q�_Ɓ�E���������mZ*����+=9[p�U��s�<��,8	k4�۷o�cr����zn������~�"0�݆=<��9Xm�c�TC�̓T;��ي`gh�l�v��IIe�o�ؾC�2�/kI�3sW��F�/RI꼴>���!���ǏV�0�&?z��p ����f7����b�
[��j&6������
�[5��1����?�5���QҔٵ��X�ʓl�l���{��K;����%0ln��r]�0lA�_�����g��aٌ�V�֋�t�������V��~�b���/Gb�0i1�xt�RUS[��~���ڬ�l��.Q�d ����2'�kP9+l6n܈�3דU��R�˿��u_�+&"ף�-�-[���5,@�N��(�޹>a�o��5;�൴�lc�L @�S�[N�:��8�EP�!,]�Y�*�@9�X}fh��~d^v�贝*�V�2DWY	fXX�_b�u �wC����]'�2�:qH�AL�(�3�ZP�xb�I�9��<�'�*��̅!�����dSC���]� t�=&&)CA�j�\]I�~6T�z�
X��(l? �x�9��8H�*y}W����}}{d��^M
	*"mx/$V������N5s��(���C?4y�oL�hvr��ց���Y:b�[�\��0$d��k���`�.�8w.���"�]���6�f#� ��򐈄���IH��g���+h[��r;%e�cmZ��%	!��X�@���9P���.����M�m��ނ����~4*<�-U��P�ņT�X�7��t�K���R�<��kc܌;����c�;��L�nX�U�	J4�dQ� eH��"9)93�"�JIr���$�Y@�9���'����ǳ�Qf����n�[]]Mـ��p�坽�0H�jۧ�=&��휁�#@
��Dn��Y[ZBq{�a�fg�w��δ&���}���a���H_��j xm���JJ��[+P���������/
�j��fh�b�U��+�*U��?v��6����+Xmym��?){�ȵ �4���F���9����U�!]R�m'T�Wl	_
&�+U��y���N|���=�9��>���f1�kN��`�����I��W/�g"�xh#c�w�H!��]��Nyyy��i{g�'x�i1 ���]oϡ^\?_%����U�N��`��j4��U���/'�:�������`Eݰ�ź!��w��gK~��y�
���b��U�����ͥh`��]��G�_�Y@��	�`�.e 5�����x�)�B�Af|�0T@�F�nA6����r�%��� :8}4a�0b �e 6|����2�I�9N��J��E_\�������|Ϯ$/J�z?�J�� ?�J�ؔ+ @ި
<�lL����뱿(a#m���[{��{���˲���v|Y�� V����Q���}o�e������ 0C�����ǏM
��d�z����g�GPكs��)����\���E�������|	�s�y{Պ]�[���Z{z�C�v>@D��eHp_mmmD�C�����w��6�MOW|/n�ng�#���y���t~��:���2������N�@R��Pel���k��iUxG�S<�q�R�2�nDd���>yBaT��:���}y��ki;�J��cכ믣��p$�S����F��Ҟ��iMM�Ʉ �9t�]iQ���:�/����uE"���*�F��0��9#��ϟ?aC@���8��g-U�'���g��:���n�I/b@� �3�:vI�[���|�UFc!lO&�����4B ��BqدJ'=���p<�1�齄�P��~�/R���{��6*q��!���
i&��%��LNN���%�7������k�G�P0�a�|��q��)P�9|������@W3���)A%j3�S�JP6��i�N��.��8�~��;^:�y^h��~��HB�C.X1�C�i�����2��� ��ځZXc�[bN�� ���).�������Tٽ� �F�JެP>���iH�����6g(������vnT�@6C��<*ג�3�E"��4�&��I�8��N���-J �rO[;rh��Zg����g�4���^}|#�q!�8\��^LB�����#�������˗�QB�'���z��Z++,�A��&�QS�_vP!+G�vg�7� B����Y�j���=z�Cv"M�VW�?"3���}6�<�/^�B	

B�70�)������(���1�����֚o���a!hX���@Y�77�T\z���M���P�1�40�	��KJbQQBX�� ������HZ���F.VQ=���.&	
</�êCR���`�=�&�}}|!�� ����|ow�9�n>��C�*4W ,���dj��&����� !�h߉������G�,L�z�v}�B�c������[)�䴰�_��a �C,,,J��-āW�+�S&�����g�߸���5�u��cx���;������
�K��q���
,�e�r�<(����.� �x=!/������~�CgExo�t�Tո. �a�0�	@�fg}�-�30R9S @�����d��)��Wƕ;�֝$um��i���W�~�������~���>�}�"d��e!�s´���yN�����e��C���$����d	`>��ɨ�Dc���}||�߁���)*I";�0�����L�"��zDRw�.G���@5@Zα������QUh���C��/�F����oW�TÎa��Xd$!�y%�H��7��6��\����G�3�s'`{Z�K	f��N�� ��}� �z��������\u_���@���<H�ˮ��㳧�����.��uN]���� D�L]خ�اpf{m���˰�"���a2hJ�ӯU숣�DY���*���,~��^XЁ`�mt���@гk����*(�OP�����yRԢ����A��'�؈���� 
��z��8���M� /��"��PƐ�l�wmmm
�hR����I)�Q:�6	DR���,m#�XwC�}Pﰋ��zK�T���sG4����5 +o:X��a{��u OJ�����G~�ػ�N�		u�·�'�В���	,G���|��
-��_ ��l�u�����P �@̀��@J�������\t2Q�@��KT\��I�b2�,�]e��wuYW��8I�!�I
��A1,,,%���7>�R��na�Y:�F�;X�E0�`T�t�
�oÛ(���;�Q��u++Y[[kf�ק�Q����y�+ѯ3Ka/bW�.gZ�S�Q�b���Y�����,L�'�n�;:����5�����_r���q����� (]J�7l���$Vo��>���y�����I1�޵vvj^؜t����Ot���#�� �!1����$$FH@X7����v��"���'`+� *-�G���F�p���Ā�-D�����6M1b�bG d���C<��M~"��b�:;;��v@�������O�āG755��O�
 t���г��wDxxZq��z-��x��ߪ}0���>,�t���Tom�Ѩ+q&M�$������9m g �O��i������;����`�C:����|
P���|"�,������ ��_�|�����ݎc=��;�מ��\ȫ��Qg)���r������+*C/���t7d[�f����>Ϥk�X��}� ���<����]:�΅Ċ
������ِ#�'��陙�1E��X��2�q\]u���=���a_��A4Z�L�F��sڀ�Nt�1���~���<z���Ψ��En�SC灷�X�~�n(
b)B༯7���:��&\:hY�br'��L��5�yp��7�8�d�m�YW`��ɴ�

bW�8�X�Zs���x������?�u*�ב�k��<��h�R3����[0٭�BAF��&lv���l��X��.�/����ܡ���˿�P�ttTo��;�@�Ng����qη��� ��� ]
<X޻��E	�_�B��+L�@��y�K��$����%�Z �28�3S]�_�*�m�;vjdh�))� .��׌<&�@���)�vD�=��_�5B�;B%�9���<�[������~yy��Q�0�.|�lO[]�\\K��\
�+��
P��a.ܵ�Z��{?�܆|�*|�
}d:溓T,�-�AA���<��OX��RIE��크`в��R���-�&��bو�l��"��V����C²xxdπ ̰l���%���f���o�����Jc�s��?c|X��������(��cA4�ar����J����M4�ml!i��mӐ§:�ٯu���H��f�='���cR���Z���.Ow��#��:�B;~�WS������f���z��nʒM2��4G7�����%n"E��yy�d�c�Q$��� �P��}��G���������y]\]��Ђ �:?�)*�8�r?a�X��<K��fWN������g����)�<�F��*ĻթBB"�pKO!��㙙��.���ʤ�e��l�i(خ�����A���ߨԹ��Լw�>i�g��C�=|�����@�{�uw�Q:'K<G��	�/� R^��F�Pc���<�y��Y+��p��3�;)��Ϥ ���3�a���H@D�	0u�:�%ȝ��,滉7ˡɍ���Ȱ���#�BK�Pp�Ѻ@� 8�<�<�Ȟ4�frE�L�{R��p�&�@ �^������n&���%�������yy��*�n�7w.8��\������6
�j����kddT�`�v��y���a@A�7�c�VVm�M�	���o��x���7�F���~� Sw��Y�%��ж7qm��y����o�r`r{�,\����%
�V����c��2�E6[O�[m�.����?p�YH��< X��pq���A:H��O��Z�es�TX?�r a��x���A-Aף�����l'�v�w.7x"""Rޛ�@����ʀ�p��n���M�_8�R���D[�4%���L?�@)�K�$bIm1�"=M�u{g^���J�&E(��L�&�l�c���*kȘ葟v���D��@��m��F�(�%xP�r?�㼿��x�/2�	#�^|��ׯ'�6��77�	Ύؼ�~�3�m�r������骓VO��)V֎��ʬ�����Ux�a�����߁�]�'�B6q��$[-()����S�������h��,�����^���<"��o�ʌ��vX�/%9��˱3@"���tD
�ɓ�F�n�TNB7t'��P��{ L��/%�Z��ߑ^�؂������] {#��^�{X��\�Fx΍��J��f;	c0��x ��?�w��ϟ�a2|��`����yҺ��84�9#C� �I��۷W���VQ��V;r�d0� �È��[c��޸��VUa�n3]���D��I������֖@/�\4�K؆�S(�6��*�x�RC^�����D1��Pɀ83b� sss�2/ ��HA�w"�L����$@
X�F�`%�K?Xa+�J�JX�C��q��DpssC�TVV�&NM�@{x�VPP|43�^2�E���\(߀j����x�a?P�0�7��W�8�q�}��Pn��Ʀp���lⱍ�? ?�`B�\o�	!�(LI���խs��%�}/;��Xܰ4���-������\�P��b�.�FTF&n�U�
�L/��^jr��6���<z(G�A<<�_�,z�%�.3J�I�P��N �:��Ba���m&҅�ZzzV$�%sP=%%��ɶ$���p�27��U��&��0Q��x��VW����B�J0�23�@TE�`{��zmw���#� ���HK�����^CJ�+&��@�wi�ۂ��iiJ�(��D^BX8�%��˙��@�7;�S��#]jZ65X Gz��w�%��2���cv�U��M���__�g��T���6�� L�?";P��` ,���G��*�i�Gڒ�����qqp?���aA�S�ɟ�
UI��XlV�Z
q��uH����g0˫o`@H/ANL��p��=�a��#(0R�ٰ�`��T@!y��L�r����|�e'�ԫof�%����,�92b<��8���1`_t��񪦦� ����^<��Z���g�����wO�k-tc�K6����LtW�q�~eK�H!x9�%w�����&Y��nOG��Ȉ��B�H��F�l�_H>�� /�+�P��Y�P2Y��E(�(:DA%��R ��Qd`߂1*� �A(��e�q��_R�!9��!}�~���0l�
�Ɇ��ۋX��.a߳I߽o ��ȭ��=��m��-S��W��[Q|(�N�Lr�����1�(K{��Z��u����4�AQ3yI�Q�j��w�H�"yS-0Z(P9ЅK�|[���A%�>����R�wkO~٣|y�l��g���Ծ���t�`Z/�cկ=��U���������W\a�<�qp��a�����Ty�ޱ��Ur����G�b^�2���ֹ��O���^	ȸR;�} �p�W�V򨯐G�
h9�wu���,�z�,p�#�+��lTu¹8��jj	&j~o��P02oi�^R�Z��չ7t)+�G���š��Ñf�:�QYu~���n�8�]3a.v�UGZ&���������k�@����*�x
}���@\��z^*_�����4*	QϠg�c�_R�X�L�85�϶,%�!P&���R8�'��u�ЫW�Ǚ�O�h�;s&?�3)�j��֫Wc����ǘ��n�_Y"٤�:�R���#�L�HY�����\T��cv`���
�:��<J�<���ϟ&���y�h����;@O�w�;���n*��JS�qF�P?ф��c5?��?J8:z�N�4b��u����N̨�JI5���G�X^e��˧񛚚�#a1�)�8VDv~h�'x���#r��<��H��NZH�pce�`�k��ꨓ�r� cɇ�L[������� 3d��y����������Ⱥ��6:!w�e?������\�+,�[��K/�~$j�pp�<�)��
@�2�cϨ�`"�Zb@��o�9jhl7�c��>�����e'� Q��������|����2ñd.@�h#�8����<~�D�Ƿ��V�5ӧ�����ob�=��{A�*��W��^�-��VTF��gs-�K@���ʩ����Hy�<�+ѝ ��e8�E6ڀ2�����N{h|zC�-��z��Pz� E-6���3b���gu�Nǰhuwz�٠)	Ơ��dm��������:j����Ð�I���U�|!�H�kR\QÔ���M'�I�d [h�P�.��"����vz��6�!:S�Xi_�N��2Ӗ��G�����[k�����ݲ���RR)�s��?W�OHX��[hτ8e����4�����r�dUWH�U�0\(l��������F�%ÖsM�x~Zz�.3�����5��"�$�5���f�\�8w�}�a'GXXY�['��ݬ.��ṈT:�[~�I����jc�qC��n�L��,���> `���[F*�TKIiEF�]��>^~��φOL�h���D���������*�2�[��7��W�5�X�K����_�N����5�f��<� l���]4�'�F�I�g�$:�4�����xԘI��]ӚuM�Q��/�a������L����������E�Dfٞ�A���堠`k` �~Nj
����^�ee�$��5�D�z4�(*!R� ws��Hw�o��C:�fGT R���������5�X4�Р��#����Q��i�j�q֥�++,��]��/�={6������rM�U�x��XD) �����LN���:�8�$[WW�"�㍬>�X*f�v�q�T�@��n�ϟ���Y�����Pє&B�nX�}kVm���XE+Go������X���V�p�邺��*-"�?Zi���y�J��d��+�x2�%��Y���X9��c ��ڣΆ��<�@��7h���\dV���7�(bN��lh_�g3����J���G�B)����J%�~�x��������sjD��+��&�c�B�ވ�$8X�^W�Cwi{xp$�֑g��`(���AQKS'#�O��^��yTuG#Ͱ�s�"���p-M�E/_�����5��ε'�YB�x>��C���|c^v��z����?)�f�!�!�o�jo@�y�0�8�bicx��e��\� U֬d�)Փ��<�P�֪�Jߒg֘kۤ�I˦�JϾ��Q��m��Y^̗�w�����/O�Dc�[��,�na��:,�C��GS����[��o��Y�;M�^��±�*�:����;c)u1_o.�1��������QQ���%Ml��/��-TU*�~.�K{n�p��ȑ�B��.��Å����,Z�u��5�.L�nIz~�h}����f�SD�u-pu���XO���ڗ�(_����pA���L�C�]l����LU+�"l��������ѓA�_���	"��#���%��2�2Ӟ�JA�t{آ��),aT/W�,�������;��
V�b��RB����Tq�F�s��{�޺.������?e�)��b�������t!�D�1P΍�*?�r�(J�,���g�Z�=�����ɺU��F�~.�p%>�J���`o��Ʈ?E�¤%�!6�@Yg�"�jx��խ�G�f���Xg���}����Q�������	�2��J���S5���~���U�%2���^�����ʛ�hS t��*�ۖ:��*��ٓ�1m{_=�\[:"��bar-��NH�����ď���"���D�d����s&ǌ�y�t���v�66H	����c��h`�m�y|�~y��ܬ�oV('A��>=���"{���ykc�fD�Lji�A�o4�c\���kn�Tт�4���M���4xs��rx�4r�Sc���Hz���!� ��]��L�C�O�^W����b��㛥O)#��Q���9ؑ��Q&�ӓ��s�bģ/��e���"ɬ�'c��m�%�a���l��wpbS��K@�&��N�gD�)�w�k���V�z�/z2l8��R��W�M.�ķ�����'	���@Ȟ��8�a3{�9��ۋ�M��S[��-�WKǵ��y�5�_���P�Zk���VYi�*��W?1f���!��*m��3�q1*_�\;�ؒEg���X�:7�q���/
sH���9ѷ�\��6V\�p��Vʪʓ}����ˏ5�i�NIW]m>�� |��� 'N����sԃ*�$N�<�=b�;nkg��x��1�<UuY�X�V����oDӏ�dwť�pڃ?Q���Z��*�4NB��=��Qǘ��4�Tš��@���4�}��H%S�l� �l��lO&���њ��	��'~s���Ri�|���C�w�37�$�C���Td\yu�_��L����$3YGL��C���� �&g>�.�����)��&��0>�(�⸓���V����XM�+�+��0���5�&����Vg>y��o��*�[k	`�=��_����W�N�,����j��O��CT\�����Mwl�=�(���%��>��I��s&&�v�I rJ��U�e�k��hT��?�(��;���n��\���6[G4���z� I��礖[��4,�[�;������<��F�&Bi�.Gww��[~����0\!�fUŃ�7v�T>2���Y}�i��G�:�}��=�P F_bT�1��+��}]�i���,:�C��]b�����c�^�^lޑ�/�.������G���l;���4xm�6��yF6�܂1�}�@��-ik)�%/ƍ�#���O��S!\��썔\�H�Z�D�wG��/ֺ�>P����Ko��"��v����z�R�ԸH��D����%R fx�x��6ְ[,����ۢGC�xA\<���[�at@A|�EEͨ���_S�@����e2���l�ӯ����;�;>��C8\��5s3� �R�!���ܜ������_���w��}�:����SL8������Ot�D ݗS�
�^��Tϰ�2�w
�9]����T;��,P�Lc����,�BV�2����I�q�իW�o+&����b�4ClR��$�"�?G҉)�{�r��{Y�o��r�������IӘ��:�Y����Ԋ����
��1��R�@,�G �tCW����Q���)��9'�e��U��F�IQ��Mܳi�wnX��P�����T7�O��؊4{��x����qn{K�J�^��y�Å45Ӯ��:]U��Eg�@'��W�e'�l��2X�i���-杙��ۂ������9���[;N�u��}�:mM�E�"�>Tz� �����PD"���S?Z]��IN�W9E7��{nn���'U�
=�i>�J�
�����2�J�&�9�'� �J��a\o��O���y5m0�&� ��7���7JJ�p|���8P=V��^z"'��п���g�`�`%�(w���%��W�/*�",�rqQ�?��z&�ag ��ͅ��k�q)'��h�µ�f�5һ��K23��u��%[������|+�5p�{Q����7d232��v�v�/���[��)/��l�잸*�βQ��31�;�@J��\�@�5���ϬՏ�5L\]v�Y��ز�9�B ���Y��7�61���D����ۭs#(���
9��S�.���.�;@�D� ^����w��=ȱ�:$w��V������R�=���hص�Z����IY� �h7-!&-�(M�(-�(M�-��&�v�/*Pb�Ґ��C�1��^/'m��Њ{Yn9�d�����LD�R��R���/���w�%���1l��2]��'Mt9��k��n;I73�2� ��/����S�\f�x��_�]�M�������ȕ�"�l�$LS����{i��ɋ"�s�;���Ҳ��m���`0����2c�(�,� `��9���-Շ���������|�+{�ό,���9���N9$㞸t-�n�,�P]�zvv���W�	f�I���蓵��)����Ӵut
�?['�yb��hh ��5ͬMcS?����͎���K>z�S4���˞z�X���p�<�w]� ��5N���/���)�8z(��1��V�b�7YY�Q�B%��ea
�uɯ�`h�	�]�CT_��~�� ��U��Ҧ^F㫘
��h�$}��V�o���Y&����=<ܒBl�h�s������jk�^X}��C��_cA0Q�gK��{���iOZ�@���}��aɖ9�^\�p�Wc�P���QVV��	->[��(�|�gB�#����	�Og�����b7�ucгL�+�9��}�)�T<��uO�bN�sB��Xl�ᯒ��/o����1%�m!��
��;��[ȸ⧶�7]51�on=ۘ����,�Jc䳛Ӭ2����z�vR'6�34�;٘ +߂?5�h�K>n)�I���U�"�ۡ������<Hy$��]�?�b�*�V��/�Ԇ�G���4���#��/�đM���$x��x� 2+e)Dqc� `�j�� e� i��o����럞dm�g��Txm5�Y8C;�/��
�fs�Ԧ���N3]v����+�|V�К��s�<1��[W)�rv|ثG�ir��<1��~?��q���z ������'&��K�H��iӎ	tN�<���C�NJ����B�#���qx�l�:���W����Qvz��}��lE�~x7��@��d����T9�R'v��5�x�ڼ��1b��sҳ{���0�SA;��ʺ�Y���o9���0�W���ӷ���w��7�-滖{e��%&�� X��"�;���<���p�g�H�v�H?�->����.�o�ɾ��xG��RrTǫ�R��`K��8��u�YI�)F�9�ff���v��������q��,�ʴ�N�D��R�qW�y���>���r;������__H3����:V��4�ބ�~���6I�dO�-2$M�����RN��.���B�U����w����'ؓ�6���Q����zZx�w!vn�*����s4�v����fD]`���ä�s��%$o��zqf�?�o�`t�n��f�̅�5�U�.H����!=5!G�"6]g�"������o������^h�{z{~T��d�����T���l��3"�/����,�#�Wz:�Cf���+ր��k�1���/�n�,,�3*�s�ڗsm�--!���U�<R�EM��Yg3��Ɲ�Vwu�\/�#��/��B�trr�'dǮ�m�/�.R1�F�b�n^,������4�v�<����8�#��x���c-�d��k�4?\ln�Fk�q���|?��{���|�������P[�2�d�s�����Ǹ�_vu��`|%��`�b|IK9�>��`̵�k�*��TM��?.��XЇ��"���±O_T\+�c=�H:�N8���o�zSN�����\e&#�����.��(oc.C�-FT!�[k�D�Q�Cu� S�>M.6�/�Nj	*)�c�y+�fљ%)+�MW�bW�f'�'Q�S5H~0�	'm�j����=��[S������l�K���mOr��ƬV�nJ�vdA$ZH���@G���T=.k�F�K\�ƻ�d%}gV�MԖ���S:Cm5�
��n=�[��9�t�SNM�gнYgf��ga:d;B�;��%���b�=,:f��T��x��1i���/�LFE��_��~������?�}`����0 ��3�v���Ng_���ם�y�ʜ�dZ��cF�r��bP�@�����@�0��~0�g�c/���h�r�̌�t;V|�o�U�uq������A�v�zc�u�4%�P�!G#��gg��d֫��"Ͱ��g
!؉�li������+���60�k�3���gy����y��`����9|�C� z,-W���W���H�I/��`;��?:n=�3�e�h�1B��z���`NY{��6�9 *��d �`�֖� �Ǜ�h�ء_]�`vL��g)��SVL������3P�.��}
�ea�A��\�j����n��`��k�J.<m�	�6������Ϩ�؃����������'{i`�����өy����;��O��k���8�s�f��8��B�$`/[� �澜C��h��+\ݮ�y�N�Rp|�����xjwt+p���W8y��O]�S_����Qv^ǣă@���<�1sU���ypg?��Nޚ��$�6{���v�9�����u�F���xI��hifZ�]dpP�n���i�1�R��G=�:N[,���β�q�����a+绛kg���Lk����<w���<cc8[��;f��g�v�8Y�.,��(&*���j�5�!�D5J�l�_�~���﹟
㓀?.���3Łu+>L��=qJ�
Ӳ�޻�?e�QL�+��a-��әҢ烵Y���v}�4�`��F'J��K�S��*����8?O��.�������2k��̺P�D̔�P~qqZ�EUb�"�I-)^YzN9�[4�Wb(Ki¼i��}����=TVt
��b�0Q��,�?��hc��\85��c�J��M�*uވ��"��h����^����� ��#ƿ�߭��0yasA?4�"��y��Lp�1�t��|�M7@.������g��#�fL��ڴV�5��
&�/6����� ����9�՞),D��#`K~nq<��N�����=�Q��r��3�cH� ��v����f�E��0����3�e��<�nK�r���|CߤO��_)7^wI�j�T޷wޑfπ	,�9���VPP�@���]W0:QIOwBE5�t�ǯg�,��?�d������Ga�����8���������j6ݸ' !l�M�'V��J'(6z#;O i���δ���q�̀��j�P���R-g��b6)nҐ�KC(�e{Պ�7��������i���L�6K��y������)�g��f�����#'̵Fa��q��@���-�P�����a���q��ȇ���u����8�T(�f4�d�h����R�vܒ	�Ɓ'}}�v���lAR�F8K�D,���ރ EuN&�4�� ��72YN�ӳ��֜�e�)+��ĝ���l��7���1�)(�7��V�}����,jy�1{����TT˂����W3�-��9TT9��D
A憘!^c�Q]����2�`RI�����F�8�s���L��x�.��";Y�;O��X�Q����t��v���'�J3�b��ơG$�ZE ���p��E����ƫ
�pٝŦ�&�z��kٚ���{3�ן{�:��n�j0<8r��}R��K�n�4�P/�Z ��yx8�D6#����3��+d��T=d�G�2���^c����8�P�u�E l+A���z�Ų5}�C]��ʋ������C=��oő]�����2���\��xЉ�f����Mb>N��P�������e�C^�|��qB�I��StH�9_��\A:.�kR��&s��0��؀���Fk+��9"ɺ =Ҽȗ�h[iy�����je_i��l�����F{�+FH�*�9��^�iŬɎA+��$�h:x'��f++��U?�v���Ii��������I���Ur"/�r��zfM'�IM4%���e��jYҷ�e�7��q%O�Ctן���%.pCr��u��>�B�� &	�T�G��P�b�iv�����\A,�l�Ȩe�n���1o��}6�$��t8[�e����{Ϣ����Izr�\/2�"�3ѷ`�'����Zv�;{����7����W+��%	>��?7Lr�X�!V��g�.k����&Cfe�v��ۮMuK\�����Uq�������?���x�B�� a�?1�T�OL!�Uo?���MTU�lA��Y0�`)ջ��ie�o�!SV���kb�H)��Qs�D����ª���kzm�_z$+I#և��W"{����� �e<3��8z�(\�:FM����Q5fvr�����QK�tA׮ )��$�c'a㙾������B��������Ѱ���M&���{|L��I N*��n��Te��@��ʄ|\��rj�y�	��;�<�]�Q�1���ǽ��JpWۻW�$NĻ�.�,��hx��Ӑhb��HGJU�*�Kkp����g\���]8�I�"��������t����y�i�ػ�J�<��y�&�!�p�*+��BF�[a�v�xz�6���/i*��Tz_�f�307�����P'�V��63�ʳy��S�Oߓ��"����#���2���kpv�3<���3�:T�x�v�JџM/����A?À`�q#�E ��T���kjY�z������jI�t�*�>\d��
I ���o�3x��_]��B]j�-��УZͽ��ٹ���,�R���]�f�=?^�`���<���ߨ̓?e)��R�''����,��u�|���
f��.;�}�_���J�VQ
��yrFT� T���͗�X_<ͶQ�oRà*���W*�w������x
�s�&��	g�M��t����;7�!�R�g1c��n����M�F�����׾&N }r���@��i
�Z�x��N{C�'1`���Ϧ�95��Hym��<p�ј��5�/>�l�R�0�3c�)ݨ�Ȍ�<�� �`�����4 nIea�?�1`VEX�ɴKL�b=�]���t{RԴ�=�r�7��V��/�#��a�?���c�`4�����ܽ8ͦ-̶U_iS��2�&�geLo�n�g��Ee�����9�0�J�&�'B{��=y���Zf
��2q@T[�Z���lR�j���;�k�ǻ�dߗ|#s)�f���ꆪ���O'�m~��Ɠ��.k�jO�)�:��������k
�P�'�G�<V�ÿ� g���y��S��SN-SK��-�@��uD�W���5Ͷ�?��FW�r�Z��� A��c�6��H�T��Mʯ�D��a������͸���)��IQv�EH�ՙ�TpZv�����[�!��7�)O��
O��ʯ��x��u־�T���`���o&����������]�b�ȵ,V��Afw�o�!�⾮W��.]�
�aQ}���(S�EQ��) 5 � �����B�մ���

��?F;�:)y�Z�֮I�Ƽ{����&�X��ĩ� 7>�Y"�k���9L |�c�	ƣ	&�)�Ƞn�������6���n�Ɇ� ��ȴy�X��V�@�Gk5�)�L�¦7ަM}�c^�b�K�4�m��)�[���B�z�TG�Z�о65-�01�����Hi&��h�a�iB��G������Ezp98r����/9t��VL�U��������*D�Дb�9��7��=��69D�g��_��)�̀-��:n�!I���B�Cj<�p���s0#��9�.
��/7�L�}��Q�M�*�G�c1�]&(�_'*����-��{NV�o�@i�QyPN��o$��ef15����ӫ�M�k�
����s�Kmg��L����!S�4����"%�ͧ$!,I�
�I����Db�ru��=���g�w@z^0]�� J����>�c�B�+�e>?ʯqFw���[�ϖ��fژ=�� >-�G��S�W��oɓ&����K�`�NX�N���zRP���9�c�J���\���>R���;-Ast����wx('��Y�;��v��}�0A�s�ӎ=�r�FJ�S1�QO�br(<�S1��ӤR3����X�[��F�[�H�X��7�r'���n��`��.iSL���r
3%���w����	u!C��m��ÿ(4������pz��0u���gJ�F����R*�M��M�x��yk�j
q�݊��h�Ĩ�qV�����^�?Z�>��5��":��,I�2�۫�w�ϾT��A'�)H <X@�%���l/۴a,�h"l�VUt�ٰ�c:�j���5�~攐�����8>��[���V���	9�W��_C�x}lz�Z�8� /��o�U5����"���j�*��	��9�����6�j3�u���UC�mZ�B�3�?�V�9�=FwH�sڋ	��`Z]����ȣ��ڱ<�lt����i_OO+��"uo!��.��Ƀm� �K8#k��f;�{s�|j}pl�sX�JOM@��v}�
7�2�������K��c�[5�)�򌧜�]�������S!~�Ie����#8�p�sUaLLL;XY�n�x�0dYC��
uo����;T�d�m��l���k3�CL�5�����Z)���.�o�k� �T/����m���2���o��]�UqUa��T(��{.KAUV�<h)�l��E9�R�{L�:O~x����A��Y���,z�Q��[As,���O�o�
1�Ƕr���W����v�>pq>���I^���uLP�}��ѵ��������[��_��|b<9�Ҹ~bSyB����t��VF�`������,��T`���r�.��igx�4I�}�SA"���$�rg�� ��yUL����7�v�M� �����S��ՅŮ��%�D��Vc7�nKS�l:�jLCD��p�t�
�hpX�J~��Ì��C����<oG���u��A��/j��'
*|��L�E�.F�JA6��f�*�.FG�~=KA����M-�L�{�h�}��/�y'��� w��|N~ /�+ϱ��	�vn�M��	��9W��mzӴR;�U�Pf�lLJf��n���H�IT�f��0c�bBb��>f)�kS�c���,�w.�U��	9�B�:�>Z��w#̀@���b�q�E�M�J]�c��l��gչ߻�[��t�xٌx�{�M<�UK(т��1���8�2��G�$�:�Zd��Iz��T�������,�#��U*+=���)�j(���]�LH�o9�0�̰��Վb���� ��A|��A��}l�*�V@ ~w-[,��tFִ?3���U�lz�����:��:������R����$����D>���zN6A]�
�^�QIЇ(Ed�Y�aRS�i���7u�ƙ�5\\Bb��?kve<�Ol#�X&�10հ���@!{�=A߬����}>�m!��H�y8}�<�G�a���	-���熛I�^�1M�-)h��-�3�-��g�5�5�O|I#)w;l�� ��?u<��,��~Ӛno��E��]���� n�g�#�WI��������Ku�
���\Ӂ��I��i�P$I��뤠��;@,���8-ױ��iJ�v�Y..n?�:��?6lo�4�e\�=�hͭӾk�'�&JU�����6����!/�q��p���,�NG)"�<��h��������#�����jfh��Jf�l*�[!|A��� �*�wS&��>����I�x���tg���f�k��w�[h !��:��O�^�9-�$7J6�O��v�E}�Bd��hB/ƇormR�F�&9�G�<c:�ri�3p}/f�4#�� i�*j]��YX}CC�Dٳ찲L�����Z ��ʽ��Z>o}�Z���orr�i�!i��\��ߘNмD������+-�: v/�m�H��!A� �X:�{�]{QF��BO���-�u����'�U����7�RVF�PC<�o��k� ��ş����Wk���D%V�2�{ Bd�I\s��R�F(�Ó[��� ����7�L�}�nq�y<|�i(�W�i��������g\�����b�+��>u�����苫r̓{�ȵp��&��� [^f��S����:��$2��F3�r攺�����}7�R��1�G�����y���������je���a��#�8(M[dv>��s���*���1���ǘ�vw�z�L��ti	�x4*�[XNc�u3�M�h�Q�f����	��;���%�o�g+Emi��H��|���J��H��p���M8���a�G�k�C�G!
�����������~���Ht{P#����V�|F���䯑�R�|��[&����%�Y�;	6��@+X	LI�� �_�c� ��j�q�qFKrP��_���g��Y�������/M�ca'K}�����u|��u63������ݯҋ����^o~v�"{p��w�ɞ`b�$���	��Y�lyt�L�Y�d=[z#]X0"�>�S(;n���a+Ol˪��=oAp?an���Wt�+���q=�b;�Э���TT8KI���Ǳ@���3v�qU�)4��o��n�c� ;��-�\�j�\��D�8}<��d_ܴEURP��\JW{�4���U��=�9_2�RK�@���������j�����ɦ���,=m#�����m��Q �3�w5�o����<q�R����Y�.�L����*v,�����h%R�a���6����Z�E7#X�mZ���.��p��Ն<�4�ns��N�!�0�M�`Z��0^�0���M�r� Q��n�������������ox��D��R�z�B��l�'�z�8�.��ND���z`{[�hoYd��
�1�=���/��:���M��R����(
��BM�D�$�%�d�5M�B�ވ�gYBeI�d�ٲ���;������3�y{�^�ܳ<��{_��)�y*B�f���K��������F�l���IIIFj�ed��߱��ח����Htkcr���X�^=�e��.|��� ϐ��e�ofX��Lz+��x�s�b݂gF�%��;<�ڵ��*׮��H���PMM�!��(J��Wod����0����o��&k�^9�?���Pc0��{<�\g�,��W��}�Ҫy�c��j�ո	�lƑZ]�u��n��Ƙҋ������>>uib�1���� |���h.ޯ���y�V�鄔#�I��r�u�᳻4D�t�T]k3;���������Θ1���v���ҥ|k������Y���u鴤۠4n���b���%����}�z�#՚����B���� [�/u�.&&&Fmd��}nӍ�T��d�l�k��4>Z�޲�%:�bb^$'>s�v~����������T�.��/�n���ԥkH�~�������d�	6�#_i-j�di�L�~���9�PR���࣫C-�&3�dŗ��Ō����Y��1���.���\�LS?�k��K٩<�N��h��z�7�Y�h��o��M\j|m"��%7��vJğ���y��Y�ً�n�)2�;��������"^7�:������g<�F�q�)~���p&�"��'�Z\��<g�6��1�l�����J9S�n�����W6�j�Ƣ�j4�_87X�LD+���tkLOO4ۅ0��y=�Z��s���t:`�m:��t||���=I�Ul���.�����_��s����ӓ�����o���ï��ދ���w0G@�.���{L��q���W�D(��=�s���/���=���];~6��N��/w��U,�n�j�d`⯕��.�Q���r�{zD�����9Y�-vx��z6 �%~aҚ��9��RJ�� _0��|+��c��]Z1#�w����5L�Xv=zd���B���k��,�v�P�Ն���v��5�w,;l7����*7#������q�y[���=����[��ol��X�����F!�4���*�OT�;����2��ܻـɩ*ߎ~�H}ˋ�]�@\J�<��·� Y��J��wzys�ߟ�ΎU�d�<rƦ�V|��]�j���dq��i�l���u#:�����M�ͫVX�V��Nc��_�����*/`��}Q~#X}��3Y��f�l n�����w]^4�o,;�`�_��6)8�:����@�L]uL�^���/Y0�J�~����y�o�bzƇ\/>��� ����=Lo��!.�=&�-�����+拄{��Wy���H�o^�`�ӿw�8~�g���6�:���/���Zt�*>�\����*�\���:rݰe�|����c�E2�j�.	H������ᙙ�/�}g�9�M�/�t��L��,�En�2���;�&!�c�3m��@�v�O��y�s\�t2�o�a�K�2no��-g~u>RNf^�������m��y~hP��������
5^�������%���/�S�%�r��mL28��-�_S�-}`5���l��\��sms���#w,��V�[V&B��Kt�Z'd�c��@QF�Pѡ���?d:�?R���Qxd>O,+��k�[L��x�8���,y�n,�h�i�!����~�����ꐐ�f�a9�n�yќ���,K6Ez���ױ[ ���
�\�xHm�Ȼ%�

���q���vC-�w�`�9�������(��)�k�~�L��|c�{g����?�׌��Ͳ�O�j/�tx�����=T�	����F-ZC�9ӆ�>���Ek��ۜ3���-�r��\߇aןM��\G��au�G�-�7��	d�ճ�ۏ#ڿ�i`zd��ЏG�wx��άʙ�'& 	��#�k=�dr<ȱܠL[�*=ykD�,�@҈۬�����~Y)W����.r�,�낶�t��8;���ZɆ�S��^[!7�'��?7ƒ��a�V�.�g����������ٺ�+mQ�v?�8�{�;��}�ï����*�X����W+3�W�i�l`z�L�S�%wy���������7:\F�rOrΙ�Y�cY]�A��%�IF3�2�i���<#/h���������Zﶁ<.�o�s�jD���SAY1;��s��f&�����"8 �&�*�8�rGw���Rg��m>=���]�-�-O]�9�x�i�SwG��ɱ��(h��p��Z��%�xf�~Y����_ڜ�·�bW|��?�<=)��]�Z[��M�,�"�BdɫrEO��aW�>�c�� ���Y�_�.��:J>��z�
g�9����tk|�my`|���\c����-��ba�M
W(ᱶr�cꔹ�7���S4��*� ��E�N1ky������O��>������0�^S��yӛ�Lҋ"_@�zmj��D����j���_[�V&���}}�.ݬ e�쥜����?��h$.��8��*���:A��;G�\�g���K1��*�U�w�o��f,~����Cf�92�-o��;�q��R���(��e{�E#�k��*�ҕN*]��t���9���,��x���&<=/O���f�]��,;�t�jHB��G��4�>m��O��"���HZ�,�]�Ƚ���v<�5##���Tt	�e�6;5^g��\��r���x���M,9�ԝ?1�w���B��H���RR܍��Xa��8�����������{m�m}`xFZ�G]�u��,�Vqu�20)�a��fYܛ��^��,���h��{F���6(���Q��rؙgZ���DH̓C�a�]�R�t˽��Ѿ߮�վ�O��E=�y�2��1���1*��:�#%�����6E=1(�$���~��ik��3�|�@� ZO��/�[�9����չ��rS)cm�J��M������i	�1j���"����of����
���14-�Ѽ����8v&?Sݚ�n�%<�\%X:@�r��X�%K ��m~Y���q�wtW����d�/p	K�i�c�4~JX]�>(d�ޝ�5�~W(L3���9�X�dĉ-��ϲ-��:9'u��p?X���Af�
I�'I�'ܷ}��(��`Luy� ��d��a���.���~4[���aE<|������I�vF�L6�:K�9��'�@�G����/8?�d��V�&S�Y��,	K��@#�4�0'��k���u�lw�	�[��}ť.s��GF�x!��S)t	;SL�V����)3�i���g���OoD�/hL'�F�p�xk~�A̯zg"����z��3*Jp
}z)��Ѣp4|�ڋK�w��S��1؜E�����`j0k��$scQ���@i�S� [y�s�1����5Y��|����(��H@����J����g�r���鐇`�bo�Q��5G���p^c�(����h� 7!�E�022�oL�����S�?5�S½�k|���i��`	��;._Xf�WVZ����+��GWY��6�B��ɓ�z������i�o����x�8�/ϼ9�}zbH����г��@�x�1Hr*2/���O��he�X�$�� �ffJ�'����h-�(���VE_���"��^É�1#S�*����>���6Z�:�.�,gn�o�g�u�(�Ýa<x���d'��lAJa:?���%���j���_ @�+�z���'�W���gn��N�(v��$��i�O��W��9���Uֱ��׵�LRz�L�SR�����u	T�-�5�w���I-�9SLФ&��l��`��_rI�4��+K�y:w����K�kρ`\i����P���p�f۹k��:��i3���"��[���W\��H$�3^Rv�Ȗ�"����&[���V��n5�
����P����m�	f,a݈!sƟ'�`���Igf<���$�"(���{m���7���[�(�4��_�c�Hd2rt��j���6����S;� ��D�H���G�=8!�+�!���)֜��Wn���J�cĥ�<���̕��x�^UUq�^� xD��cl�����r��>�����[�)�;Z�}�m5l��x��]�:\m����|���z���H8�OE��������O��n	�~m���	r7�E��5�>&Wc�L���JR�n��rc�W���u��6�/6��С��ڨ�3�;@���#��2Ĉ�A�J�I�ٶ�6���aT�UU#����r�>�sދ�	��vt�~UQ�v�A��?���Ul�qLi��6h��[�Hv('���%�_A%	��Vy�:!��[� qT��ы�E��8�%XE8 �E�;���Ȅ�Waҿδ��;��cvf&�_�H����K����;R���V�6y�NOѵ�Zl��{�Nl@��u"ٸ��U��샲;��o��hGx7NRU��V�P�HB�]��Q��Z/��Rp��Ԏ���{r�W��㾭���Ub�B&���H�!�����_��Fw���t��!��l�)�+�rg��R�����)ہ<</�p�ۅ���o��*�L_t<���"nU���#I���w��� �(� l�����@_�~Y�y����Zp���Lk�S��Q]>���=�8��~�צ�U��ik{@&:��x�h��'�����=Z.E!�~Հ��3�[	��x� �$��0��e{����P��ޏ��'�g�5R{΢��V����8�
�=0�E�:u��X{$Q�b�^���S�!a�t���n9�k��s8�NP��lB�p"�3� 8�̔�llB��B�h_'��IZ�+�dZ�a�NB���-��h��.nt����{�����"�:�Y%�8���0�]`�/���5������{�?��)W��g�h�b�ȕ���@�h���p�u� qm�W�Q�b���;�	&�?��J1�P�+5�YMU���5���OJ�m��Tay���������m��<M{oJ^?��$��t�%�@:ݛ.eG�|u�CT[8T-��9������<�.���T~tو�3Me��:�8��G���i��`����w�m��٠�>A_����R	W���&8��Q�eM�� ��γ�u����U@9��u�ƛ_�hf�*#�����h<�	@%�*!7��-�d=������T��?�Q�6����n��qzfB\��W��D�N��"�}ޱT$���s����bBP�UK �����.35�`�dީr��w��h2����EP�?�_ߘ�W!�,�5!B9l�ξ둹��E��9�9_z�l��@}���y�C*3��Ӆ�ڇ�/�L��#]����[�NAݺڢr�=�����7�;��`��Rs=;�H�4� k�z�E�U���x&a�G4�j{~�5�==���J��?	�����q�P��\ߦs~��v�C�&%&�'�~n�*�C��S*k��uN�[iЊ���AO4����H7`cERCُ��It����o���j�����q��\��G��FiA�
��p��({�0�l�ך��@�d9�j�
fH���]b�l˥48�;�]Q�u�ŏjG�ȷ�ŏ,;?�$|湚?�y)�A� �|P���"_�7�Wy��W�@{�[1=7=���+�B_�k�l/ ��Ϳ�*<uҪ�#}��Z����R�x)��E�yL,�Dx��g #(V��h�������T����6XHc�~�S��	@j�:,���/J����E?;Ĝ��;>}S�:ؔ��+�
F��rJ��S����k�i�����m�W�_��lGF1]����o	�.eR��">�������]���� y}H�
Ņt��wKx���{�Hl��Z^�K�I�S��i����*�L��@�5�ހcV.8�&>���E���;���ہ ���*T5�	�-z�`l���Q\N�7�n�Lz�����@����,L��Y]�:M_��2�y&�b�a�b�ؤ*7��${6��X!�^��\�H�����"\+:���m��f�n�sl�L]��F�� 1-?֋��xl7A���ȳi����J^5�� ����$��U$C?�r�w�oL" ��Vޑ�C�m�Q���t��_���`��YH�AM���H['ʥ��lX&��x���Rrc�|��@�Q�m�j_I��أY���B�= ��+�w����7����e��}}�~U���F���4���l�4�@z,̰�g����H�17�R�_��U�Y],�9k�Fi���JΎ(�^����#\뎊�B&U*@�M��O��[��̄#�*|����ͱ�1f)$�}8K�J��U~�5¡1�o��^���;��;�@����_r36��ƬAA��l�e�2,1�K	2���C�%LuY�7Z� �]J(��d%ˑ�PRV���}5>�"dJ��"<#H����WD����b�W�M�&vkm�g�+�L�2�T-;��5q&���N��D3��vg�T����aP����bc���0_oU�cD��j��D�qe�v�N�2���n��/���V3�HG�����f]�v虜�,2R�g�!�'@KE/�?Z�B ،�<�&�ylT�i�t9�=�it�cEe�(�ȭ�$ mF��졄P�[5�gF�a'�Z�q��Y�ϳ�5�o_��ӥ0}�Ɂ\�1��, Zb� �dL������*�4drCqZ��w�[?"�����.���j��'ٔ�h4�����Gp�ȳ��[t���'>�g�����魮A�L����x��=�҂�1z�ǳ��{7�� T�,D$md;/2?�]��w�ژ9D�����觗��l�gtt�x������-�>'((�$���n$�ð�"�(�]���{��0߻ʂ������[�g6e���ת��&T��Q��`�8�[e	�%,�+��񾺎�hu����Hv/qP�£�|�
�C�M%��[��.���^6������Ծ������QA�!8`���?P�ʑҲ��y�Unʙ6/-/�(w��$K��G3�٨���w�v��I̔MV$ e�0�H'%�L��s!�$���%ؓP"MsZ�^�ƨ�\�G��1�"���R��BUI�V����XO%��r!�4�lݿ	'L�����_���/���d%<ܞo=8�y�+���D���񮝩�+L������Q�ǳ7��`���v{�`S�x8K����I��@��4@�r�k*�D>��|KX�fV]p?���6(� V�T�w��M�CI&� �Yv�-�,����i�.�<XS+�Q�* j�D�8�G6[�����L�"~�pZ�`f��{RSf�+N|`Ү�W߀O�(�%)k��[ۃg�6�\gF�@/B��̞n�,!|�6�����%ȱ?���Q[k���i�T���������>����� Ly�X����"�^��R���k\{ .���� ɝ4�B��&>���}⸼�/4v�DF�����QZ�5`�r�� �#�;e,�� 
��'jD֗�O��Db���*X!{�hL��bv��X�RŹB~�B��2?񐔼-1O�'Yf�B{������0�;g0q���wl`r��D��;�l?�b���Ͷ�����,vV��9��\<��r��-��R��د�qߩP��j���O���>�/�1�,Ј�M�&� )�)�ǧ���ԏ��4���j���h,P�O;�X�wy	Pu$Yu��ʿ�Q����=;F��WWO\O��y?���v�$ڦ:226V7��F�Ȁ�l7�fLd"�r�H�ҽw���m���-�6���{ ,��jv$1\�FZ���
`��Ϳ�sIX	*�8��s�˖�N0��ig�D�ς����\MT ]�nÚ�x��v�anO�����ݿ�x�>�T�X1�@��'\_2��\tצ-���Hd���h����喽_^��Lu�����͚���0\J��~�9���7��&�:g��S���3fgj|�fNA�]/��q��{�'lv,t*V&X���߿�hI�w�_��la�U�����#��6��${�f4�&dZZ	�'`�N����1l�����"�J��!E�|�5��FFۑ��'�`ɀ��Z���4jPfo����]�g����������b�5��B��5b����[R'GM�x���R����&�0�x.���h¼U�?K��^�>�E��އHzh�#_�Ep}��p�6�}�S��I�N���߭�&�������8�L��uI�a�5M��~5��9.$W�w�-�Z�t�(���4P��·���' #mu~� ��s�]�$/.Kފ���W��qS������Y1�!�8��W�v�z׀j.y�y��W�g� �n�i��Ͳ���V�x��=3{�G�ǰEZ��0��l0�jȰ2�Նr��2R_=R��������@c���f���ysm3*;�w�災%�on��*\nPF�^��]��O�" S!#��8�h���:w�bx�
i�_��]N��	��/yksrb�%�	����q��
~{Q����Q���ݐAmX�a��?~v�`�L��wF Q�}��A£���;��g��6��A�Y%��e�p�Q����k;�$a0ʢ:01��`}���b�ױ��Ó��~��@���K�$Vs���>8X��M�X�&ڋ�LOx��ȝ�O%3c�}�-��I@�S�bWFt"(�e{o"������LKpYٟt�X��T��ǋ�~�[�ل|����+����3����U��"����>V��G�K6�)H��h�q#��8���l��ɩ���*�}:�l�dD[v~f�hm�au�{�vG7���dS�b�׷N���k�P�xı��r�tjD���>��G@���˷B�^��2�F�Ǔx����+����� 7�7V�٫f�y�@�h��/!�8�;Q�}��?/�X&�6���>߬��Q�#h{���>�wWߊ7a��ގ�rTL�@@}`����4Ǔ��I��:v�=�n^@*K��*!`̸���+xӪ����b\�M��	���x�>rc����F �#E�6:	vg��DLKV* ����+:W��vI!ԏ��kWi�o9�C0<���{��BB;o�:��O&C��9�홹|��k���զ7�3��b�V4g�	�v0�(�j��OQ�ݡt�+1t3��$D����h���� ��8��)�tVhcϥK�?ho���≶nUU�p"�F��k,	+q�n�z��:��{���mb���5�f����q�Ӡ��h���������Z�����,�h��%#���l���!_/p~_b��j}�Q9ܮ����s���)�� �u����י�rX���)�����ҟ�?J�Y��0)����<3理u�I�^ml���y��^��n���'ˎ�6�3��8=��P	_�f�XrR0��$�}"%k1��42ĕ�n�	w��dA]�Jc�_�P*��3�� x����'G�8�x
�}rrC����Vt%e�
a8�r�i7�`��+�-Y��(©49:�gK�ݐ�,Xn�8���R^&�lQ��.c�<�7l�28�6�C�O���| 4
��������;��
������4)��:DM6�n��z)�A>� �#bv:��ΚQA���eE�!ޗ�AK��$�����i��B����eSު��''>����e�Lj%�?�A���:���Ew��/���Q���]����� �<rɖ&�& x��ߚ���b�;����Xa��ܛ%
sB=�,:���ju|� ��Y7�:��-�9\��#�2Y�J�o�@��$kT�����������y���7�$~�jH���&��F4�_v%`����I��`JFת��T-�਄�9I҅����!��'�m���ī�)(y4@��pV��vk����/U.��;��7��-L�s������p���C�E�W��Ԑ|��F��QDF���"�����H"�w؛�M���Xh��Q�/�?���e�t��8�F,h�����"7c2��"Kִɡ@=;����� ���@��t�4�mw=�r��1�V���d\���c$��L���dg	p��_?Y1,s4w��7ٍ�\���g�Bo�-5c�nr��΃(��i�fɺ��WTdj;��L���*����ȳ�+�3	&d�SOȷb��4�}B�j!;�]ƨd���e�,�y�2Nd3S��.�9��_�:�ʖcg�-�W�{�#6�3!6���ur3Çѷ��y���FJ�`͗k+�i��z�x(9��qW72V�n.J�}�1�#�&������g����1�p��
�i��H��¡\~ҵ'^S9#/�Ӝܯ�8���Oӿ���ʳ0w�Tl���Ti���������w-�¼����MR*w��H���y��Po���V�&�^�kK!��j�h��-���&�^��N����k��[g�E���sPb)��,�!^���A�O%������g)������!%�󀾴�����VPk�?_���I֖˹m,))i�>��,�טq״I����;���+�-U�;�OC=�t���|�O�z,�Aޓ�3�$�_��kW���S�]f��?�Ĉ�(൏�����8�\��bdo4vC��H��f���7��gR��o���7$�O��T�S��9��!�!H�ɯ��~����v�7}��p�͙V�*3@�`���8CJW$���oN��m��r�{�*����ߓ���P��<�h�� ���N"o;΅h�{�9��477�
��O���H�N�A��oM��2�ID=���/L�������`@vٮ|g"z���ޚ�wDfw��;V^��8��< �q���@���X��ޞ�����󘗒c�~_D>0b ʕ��P�O"55��q�(=nj Ge�v1��t"�Y���TV~�y	����
��X����vv)0�H��.!�Y��[�J��ّ�o޸ͻ�m��W���226
��J
`L��H-?2�-��� �$�n�F���?6��{��ڜcֿ���ݫ"��k�Y��ח���c��">�o.a�74܆����G�*^���FI�: ���I� ���)�%*z����[�zb��yLv��q)�.��sr�ڣ����D�u]��\���� ��<J齜�U���V���hs[f}�S[[[�{f�J �"�,.Xs��tP\e��5R��^7���"bsy��%��.bN��"pd��hV�����;��d����\܀�v���d4A��\�J���߂�JC�#êƜ��j��o��CKpA��I�(�����a� �u�z�߮�R$���2�,���U��oP�%8��(�.�@n(?�_lS�B6r2d����J|@?X�g�y���!:E5I/�� c��U���^5fFĻY{e���'��?7Jۯ�r�
���+�PA$��B1G�t�Z��=/�S�m/���{����jO��%��M���9�v����7�V��N[�����f�I፲�ļ�dS�ɕ+��������G��bY�njnQa��i.�B78�����O���24���8 !VSB����Q&����?���^ݭ���������G�mNڼ9�<@q&$|A�J���mYK3.���TRo�A�{Kwi�4���˕��mETVH5pV7UE�v�ӥ�¤P���T��\�Uf��nl4E��'�,��B�e�wY��L^B�f�P��+�}�w����iR4��^^�輯��<�|�B��.X�a��`sI����D��Ŭ �$���5�q�N���0�)����ɒs�yO9lώ�S���h���Yy9Pk��~qq43�n�a9Dd��?L���.3C.���ޅ^E������/���b:�ҰD�&��������骷O{�(�w���r��9�N?�}��UܫI̲� �
$8�S���`�KēiNc#��gW�~l̲ѿ��H%����)����V�U3��?����7_��M�HT��7ֽ��h��W�:��~�|-���w+.:�N��O<5�%�<�j�'(p��`�/�����,�q2Z�8S�,$u������ �I��ԯ6 �#�#�EV7{����o(=ۀvI�u�O���q� Xs�~Ă����MDN3�Ej�Z7]	b����`�����$H:�.�m�?!qC�LU�[��H��MQ˿#�nZ����'ݎ��+���e������u��7�W
�"��W-,�L򐘄]SK��ۇ;��:Y`锛F노�k���v��n���	b���ݗ����S�6x�V����O$���ĸ���W/���7,_��yq����TF��TK���M5�����R!{�x������i�O&�𦬉��㛳��E����������?-���D�����q�m˺p	`�.I�ɑ����4���O�$��o~�y	��9r���N��`5^��Ϳ�#ֿBk������G<d�dj����$�;*�M������	o��^��sϼ��-č�m�ߌxn �� }�4��l����&E�ͥ塷k���E~)ѮTE��/��F�'�m���PT���l�m=��WC?T�Q�ڞ�C�h�m)p;|�`\t�T�����aH�# l�"�%cA�w��N��K��r�|[@����Y�C:��f�L����$y��6�^.o2��JUZx�S{�����C%TU'��&�+G!��VS&MPoZ��� 
�4�{���W�w���j�i%)�m�#�����ߜ��ͣ����>��i�K{B~ۆ G�� ���`'��*�&��'��z��ojྸ��K$=�d����V�5YY@��5 |�=4L6pPI��Iqߍ2^0̮�˨��F�],�k���	U2����WJ���`�ɂA9Ř��jr�P�y]'7��wHu��^R"5��8�ZJAW.�2#��ܣ��>]����RO�-r�|���פ^L��cCN,qj�A��7200 �ٵG岓i��Q�e���l�55�G��t8��&�T,D�?!�FF��6�;�&�#�� ���*�B� B= P0 �()R���H:ե�Y��oA�bV���Ѐ��/��h*�5y-"�qy���f�������*��w�+�=�a�v33�|�7�8�bU?��n� o	�~p�V�y�\d���/8����V��g��8�R2�
��W��*5�u"�e%yCs�!�-���F'\��{�W��=�Ž��o^�jr�.��`�uC<O�wc��:(���$��W���U��9�J�#��i�Zd\g$6�8f����R "�n}�p�.Pq�BR3�B"�Xl!d%�U�[�~O��_��Dk�Ϟ�*��s�X5�Z���8Gf����UBos)�Y}``���h�w�С'�b�E.a�L�d*ں�����_7��}��K����m�l/o�$�
��!���_��˯��R��>e�{��Y�nK9���P�n���n0��0�5!��7��撥�GX�h��t痜���ז@�rO� ��ᷚ"*'��[:2�!�u�y�))�!�(�=��Bj���s�.���k+q�k���� W��D�B9ڏ��O{�G��'����ɇ�6�?�����_d� �&���wE���,)�s9(X�PbU���dvR��˹�R7���w����0@7p[�ՕS1��:IW�e���L���_�P��迅��%O � �Y��P7I`0��7��C��'�.L��� ��Y�����ߠAю�u~�e�m��M$�]���V+�{L��1�o��M�/���������I��J ��з��wp��G�ӟN��i+�c)��C1�����?
��.���n)Sb36ұ EYL�^�7��u���?}:Ff���������ƌ�wEՙ�'�Bĵ�dv�Q����0���CAU���V:뭔-�L1}��su����7�����#��d�RX��a���^���u�A�~���n�Ŀ�`�6T�C`����#����`�r"23�M
?4!�=�O�p�dē"�e+�z��'kNZҕ������m�Ů�O�\� �i#�%��J��M�_����ad/�/������,*>�$���
�-n]@�klj����o���?�n���<���c�k^����}��������{�D�/��>���0�0�<��Ҵ��<�Y`z�+*�=9���nAA��p�7-+)<�>����ĸ"�L�K_5��Q.�@��vu���+5�g���o�e��i�#e���L ����V��|� �F��Q?.��4G/IH����J�%`&ޕ�����'�%��3)���t1/��4������ȇݿJ���T?��+܅�#��Z-A��3��q		H��G�,���!�\���ᦅGA��t|w��Ne6�E�#�S�z��lFvxz�rH!R,b�n�J�H�hf7]�i��d�zۡ�1")�֟��F��`R��X-��Q�W�^i�96��<�Y:1{B�p�`�_��@ 봵�?� 2����sӹ�R��F���y�/"Т'����s��HGQRNN0z�eZL��'�����P�����wzI%�Ԭ_C����)��g�|A�ս,�p�	�|>إ����>5��6�ih�i�ȍ�Nb���n��.痳�hnn�m٤�IMJMe�|����&�O������(ĸ���V�K��<}0�h_�sG�z��Y���;�|\\d�u��;@&,W<ȢY��m��#�����9O ����C�����(=��j!*7o*荎gڔ�e�1=D�����^��[�O��-]�M�s�&TKa�[�w�$����7cy��2�A�ڙ֯4����u���~'�`�����7D@=��Ө�t0� ����P���Sdg?�d�02�H:��

�r�����rvW� �ǜ��APxT ��N0�a�y���HQM�Yvdڷ�����.W��ICCܖ�fm*�RK5��4�H��漉0b\��P.�l�/�g�� _ so�~͵��2���h!(��X|��$f٧������һ�ZSSC �"�j��>k���E��Dz�5t�K�8���z�!9i��+W};��Y���L^�3.�K��X�*��z����dɞ�lK����2�s�W���ՠ� �ǅ�Ї��%��Y��B����aoQsy�P��c������E`����|X��S�fޅ�]SM:�n�QϾ�� Ϯ*a<��H-����������@����,�i��v1{��Z��&���������OB�%V
�:�������8�i�Y��e��`J_��|��[v���|�P;��ʧ�Y��O�.��jS��UVH��]�1<p$�g�QdA�7$n|xq����}T�o5�����"	�?57���'��k��Z�B��Zʵ��"UI��|)~�Cސ�2ˢ;�=��ב����*��r8�3�s�,Al��2��$xv��-�YK�6/)!| n;y;���`SF���!y�3蹞�����FQ�o�P�Z$%'?D��c���p�#�|�[�,�i8��,�Z��C��]x0{��؛���'����8��3�2�!*+�V�H�
�wu�.��!T��A���Ch:_�|������7�C�v�X4����)o�p�ᶃ���k�"#)M�HH�2���"�V	�1��!����q��:(x��z�|k�͟�S}	���&��"�z�1p���������B�
�q%�/&������}���t?�	�v9]�Q�|7���F6���@A5Nn�O�D�_^|���}�z����+��GG;|� r/ bYA}�t���d�������>�k���B��L�������/�k-_w{I�b���l=�nC
�i��h8�VVE_䗺��qj��U��'|�ȑD���ux��XB���) �]�%��Q'�h߃"�ׅ��F��H<y!�vI��j����M����A.y�g�ΛU�s�A�[j�"O��Q��b�Ή�2���i��°�u��KTBߗ����B�?����Oɸo�Ƚ�����*�]15&�I�za���p��@\U������#�WY)U9VC*�M�!=���W0UF�Dxu}]
���C�\ޭ7ZJ��[��xIÆ@l"A�*k�B�c��M|FRe=be�&��Jo��'��J^J1���9S>�* u��X�+$}����9���J&7;�}<�����Ѳ��//��#���V��m�=ڍ ���\�eQz�c [x��~kaCe)E���j�ܢR�jx1��9�Gn�o���n�!�p��?�B�W,���D�j��o4��8�]=�?_��p��,�̄�D�dxbL�}��� r�%r7rBFi���2�YP�4\��%++x�3�b�o�k�vus�H�#���B�x�1���	YY��eDR*܉���w���:�_hΰ�GL�K:72!������o��7�4E��]�/N~�8�� ��.�_�?��z�1E�)Ù�_��{dg����ri��[%LŽ$��P�a�afH@�����X�s��"7<-y"T�����J��a6⸡��۬u,�C�A������#���O�<!))k���a�4�-0�L��T^�F$���"I��t��n��C�C��1 ��>{���|+^�Hm���,�@��Һ�V��z��߆v8<��Saɢ ��̃3*g��Y��@"l�Fi����𸝧,nuSs��G�e�I���`�,�Q���A����!����[(A�ȕX��H��Wx�Ȋ'!Qkq����;Hf]�	2 D��n~n2K����+.Pg�XЉ����T !d;
\��7��[:耾���
�G���R�9b�Z��smz����|6/����Ka���R���Y �� XX8�J��� ��ꅈy�u���}���	%�6�
�x`�Ӱ���E-Û�Z�{����;(I|��yU�N��5���i.��h�r�|9p+�'v���ֵ]L%Ԟ��3�įh41c�h TIii�PO����h�$����7ϳI��WAꕺ0�&C���>R��F��R,�9U�:i�^߿�M���g?E絿���w��#��E4yoģD!\7]�T7�-�<�(�1�=0���ȍ-(.���'�4֣ffa����������>0G�'K<`�(G-P�(���E}"Y�������V\*������.e�r��T�y�H�Ql�Ic	��V��i�(WF޻���=��Z�����[�y��H���D<iY�$kѾl�c�j�ȯ@E��?����^s��W��_�R�>�Y�eW(�J���%���d�QO;���������Oi�s�Ο��ӱ���L}dS�a��WHGd)F���+��䑂R��ʫ�FD�� �*��K;��@�8��la���hl��KUB���O%P��V��͸)x!ǻ/��4�r�"�pƦ��V��g� ��sɹ��ȕiA�W���;����R���w�.��ޢ%��Vi�.� �b3<S��')�����=^w|?�Cb�(�x��qL���4��4YZ�A-vv� ���)d}K0"
��t��i+�ۃ'�gsgQ���=��4]��+m*De�AU�T�7��e�.��р\��ٹu�h���G�F27���]��g��O|k�v��a~�[`�۳7A'�����k̀���-o1��21hǔ��x2/�t:C	�iR�G� 4����hL��p�M%���Ӏ��� �2.fq��ݶf��E�Dq]V�Q���q���dhE��Wl�hW��u9T�"#f�/�$ͨC�I�˴�(�n\�ع�Np:�2��fͱ��k��b��6��D����gb�h4���L�{om����2���|~}�q�yn%��rJ���

�_q�U<�s�rh��ܙ�������]�����w�"2�2O�"�o$��(J���"w�8rQ�����^��<=� ��o��r�P�҉FF���\1T"�-/���Y\r$[�v�U��+�-��oi���͗��+�,n�}Ob����h��k�Rpe�8-=݀Z�q�"ДJpX��zKҖ�Lk�

	aK�
�]�����M��E���?�+!|��Q�������z:�>\C	a��|����F�1\�[� �ߌ��\q�F�f���`�����M�	B���ke�n���j�����QJ�ѩ������Q'��zd���C`��c_+M��k�O�]����9��l�'�h�����|�s�q�k,�RO}I5gW1�QP���ƥ��Ƥ�T,(�0K�"!ʗY���uu"{���dn�d.�/|@t,\��.���
��w�gv���"�:"am˯��Q�u얯��Ă��7-y�Ѯ��4�|:��k׊�^9T��M[��9�9�h��]���<����k�VE�.��V_k�w=���s��"m��C�i�i_�o��2S�IS����י���Ɵԡ�_��V�H��5��ٰ%��n�ꥯ�Z3Y��ьށ����\��(Ϸ����f*��[���n�3'hY�����QVsD�);�M��f�<����t�2i}�4�Gr��#+f*�gT�Qc&��*?

��Xrl�%Mg����ʽ�c�,�t.4����5���� k���M�]����ў-��+;�k���g����:�}���4$7�[)��P���:��{�T�`2T{a��O�1T�x�4N��fY̩��֦��ϼ��^%�E���������<k�cF0_��A2�C89�ɉ�y���-l�ظN��1.�olnv���k��U�&�Fh�Z��`R!g���Y���`��l뼷�Γ�Ƭ6<:u��b���sJ;��=6�p%�_L۴��=�Wzyv���0:���H#bܑ���&Vֹ��4d�>E�?c�/(��DB�x/��ʽ%7|1M��&O-�U8�ƲV�A��'���&��7���ivx�Ѕ�{ 3��[�Oen���1I��'K����HK+��QUn]�]�,$���?��7E�y`���7�,����J��~�t����������͍��ŗ2��1���y����u�FC1�:�{����'��c���~5�?l*�9��!�DpL�W/)�|�N����`��Gw-Q�f�T�o$�w��ѐ
�ӧ+-���Hs�!����0���E���󎮏#�feeᇉ�`����NN�-g�]�VW?����u	�������j��0s�Cn���V�	zY�,�ޒ������3t�#�_������,݄f}������~�s������c��/:Z���y�r(��������:{����T��|��k�!&f�Ċ������m��V�~�-���.��)�U�=>u�DՋ;w� �T�F�� ��
�sL��$�흛����������oު�;�󥵛��ieF)D�8ў�'B�`��T�8/����XzP	��8����6��h�2�58u��2�
=������ݼ�u��^N���i=��w���� !�#TN�k��:ȆD��,�����MT�"T�k݄p�Uf;�X��Py�YȐE�)���(���<M��R����'-�`2 0���`��J^2Z�N֒����鹭`��W���o���X-��
!%�!**b}j�f�J36O�ut���Y��T���7p���Z��\�7���;uu�<�ǘ�>�}�"��d4$�y����[H�Q���P��ezkh��h�1��u�\��M�e��2+�Q'`�rL%7��[l��'Y�=���wp� �n̞h^����G�u�Eut��F1*c�H1�(E�� �(J�"�� RX�^ņR54�Ra�.E�^E`i"�KY`)��ܻ��|���{����w�̝)�cd��W3=�f \����JR@��F��Vr{ �ˏޞȃ�F|�_m���qZ�V�SQ�:�`L6�37ڂ���w�%u��뭇���Y��.'�bHv�-at����U��nw�W|���nrQ6)!b����ݽ�y�J"�5��&;8}����Q��P��4��Z��1Gu��9< �9� �W�c���!�D�b,A�} �b����4���].-e��-LO��0�vZ#� �o#))��2�z>�]�\K
���r� /��Wc��m7�+q�"�wpvfL�y�U؏"x�zl3ei�ee���;F[�U�U�����|��i���R{�������NAy�#OMo�����5�R,N�xX��$�^�֫>kщ���Q�Ϋ4����@T>� �Vr	�{2匈j|I R��4�r@�EH�5p;�_��
($17�nw���9�-�Dj{�~c�_��ɖM0P�ج�f��)���nt�R��y:��]s@(dW�>ή��w�}i���.*��'�F\T�j/�z�Nl�,���ܐ�+� ��	I�{�\2
��&g���0u}lsn��T�e���js���>׶?�M��[�D��8p�;�����z͸o������&��� �* [�u��7�5���9-퍁�%�SQ�DH��'��)==�x&N���:18�ޓ���ڶ�ኇ�G(����ӊ�w���������U�M~<6�ڍcQo:' �n���a�0F�6�\�;^N)7i���a�M��!�:�5����/	L:4���~���X�<�_{�-h�;�h�z�`�l��ԥ�ը�����%,�W�?��Q�cSdH�}z ��=@A�[��ňX[����S�p&"Q7+�
p�����I��Q�Z�D���xZi_�z~��%��� w<(^^�i��Fx��J  8"�f $��,��'S�ǪD���j��d`���֯�	��b�Q���0�P��?� �J�H&�E�쎂��j�_&�Ey�F���"m�ѡ=/���2�y��\.�I�#60��̏c�G2���.yt����E,�� ��(d�j
8��#�p�D16���G����`����ޱ��GL�v�W���DTk�9����?Ⱥ����1P�S/����Ťo��2�5�Y?t��x��~�mX:/�U�=x�69Jb�\�$N%�
Ċ�(B�c�4S���C���G�����l���v*Tq��T	x�*V��{�J�	�0���L�f �=T��,__|� ����,���q#v��ΐ˟^¾�on�; =
��<^Ŷ��Ch�@M:<+��*䊠��[Qa�����%�*�'�;`܌�B�ؐ��6���]t��ki�;H�9�9���z,��a�@����^���z��~z�	_P^�t^d�F t!߸����3~t ��rS���['g�V>��hv*D��BPO})t�J�m��s�P%r�(�x� -�� ��N(ŏ��q��}2+�v��%B�BK�����@X��|��?��_�K��p�%(��=�
�D/3U�h(؀�Pmv�3 :��F.@��G�s�-t�ŵ��ʵ�/0�����y� .xTe'�},e"aw�	�������������6������.��vV���!�4�L[�L�a�!��&O�nG/6�<0:���g���f�}�<��z9yoZ�2nk��F�+a|w8~G6�c6)�G�u�<�"˲�0�QQP3W\�k\N��+l��9�r�؛JK�GOgI6�F$�!�E�(���w�ϖ�2��>�� ¾�R�7��!Z���xb���*��J���HN�C�m��=4�����E>���NA>�y�MXo������ �BP7^�>~����'pѝ�6�����]]	�:k�kH�P�J�zO`�=��q�zry�����6��!��S��Z��GN�����m���D�ku�L{S�$��S�v�`8g;�1��A�7�zR�Q퓟;�����O���Kn8!�d3��E��^���s*o��������`Q�`@��G���C������#W|
85��OZ��P|4�
�c���rP��S[ےl��h=M����z.�q[� RֺT��m�o;o��F�ah0_���A��oT�:w�X[F��3o��AD��7Xz%�7
��6$�=5�R�^d ׎E���9���+q~tC��$Du�E0��
��Զ�����Ц8ަ��oTP��|�M@�D�^��CN�����5��M�w]� 2�`�g��x��ax����(�)�$�����_� �م������{�aVݾ���&�9x�"P�	��S:��VOp8�̃����WIT��C�˲yqd�Q����\^7e�H�E��[ͬ@���ӥ���wN�3�;A�c6���mb*�۔TO�@ �������}^�fSU�LDe�cy����={G,�� ��c����I� �[r�1�n��9Iϰx����*�8�]��.�q]�	�|xR�c\��A�3��׬���2���V�N>�F?#���c�06��!��j�����c�ZA��{�G��!ѐ/Ҡc$���U��m,4
�����=�¿�h��34!�"��'��P�P���e���#������������q�$�W�2�.^�:��	ňXR������f���^�[*#�����	S�� &)2���/ρxF1��F�� ~�M7�Gg��n��x�mj���&"�sbGs�}����*���߶M�%,z7��5�)�W1�X�>]d�3�.���Q=%?�J�; ��p�"�[�\|Z�p��#�F�l'�+����xӥD�r�@��S!��A���]��czR��DJoQ���َGٸ=[����|ja�-�C��D��� ���W"�3�2:�5��c��3$ :=á�j�� �3��Մ�g��@���b(�LԶ�<=����ٸ�%�Bȓ��[�tZ��&�*���DoonN�}��b��!)���c�� �6���0|�����V,�O[G���X�}�Y�S�b��	���{7�6�Ю�8�cF����»�l,ԍ���t?`v�����G�'�A���Ui���e,��`*\E��<�@��/�;>j�PN,�4~H�SV����dC>}�]B �M��R�Wru�	x\�Z�Z�F�@��c%�E�UP~��F�a��:�����Uos� �P-? C��S~�C��l\�(�h�y�ײC |Oڱ���mA�n���x�>&����%�y@�Y��}	��A=݌����a��9n�����'�'�6�i�&2�����V����47�l���a5�̈́��D�;��#�����y�I]6Ρ��$�����F����x!��w���S���0�4������)�/�qd�N�FJ_� ހ���s�m���XL{� cZ�qy�+�/�"�VJ��}s����MT/���	��v�4
1�q5��t�8��vOJ��~��Y$*&5��A8��I����P�������)}��j|�[��ST�ȿ� ��D�@[hQ�� �c
(~Xh��&? �M�?�$C�!����&ئ-�혗(���V�r�j]��\๼��Z����Y�,�B�6�!T�Wb�~�8Gao�n2Aױ�ǧ$��ۭ����Ș�/���n�-cv8�s�h��J�����������Rj�l��C��/*���>�;ji�j�>����I��M (*n�+/��GV�����^���.��5v������^f_��A`x�G�%[��v��=�Ї�1|[bX10�.�ur�Z
rJ` �ʫX��K��������i�8�rA�: C'��D���*RT2�#��kk;�\��ޜ\-������U1�'8m�����ѨY3���}rH&�N@&Ƹd����`NW*>P�'��$
e�urU��mRz�t��:u��C*F��a<���s��m�:��#z	�^b :#���dol��h	����:8����~�J����a0��V9]�+��2y�4#�Ţ,��Y�$��[A���	�Z�����4a���kA�������B���33ڮ��/��"�h+Ȭ4��w��W��x�mwP�v�|�'��a��f����BxU��p+��NN	�d����Fp{X��)�����q4�bbx��~(�����P~,74�Ȓ�"�q-�r(�z�r�OS9��h]J����g�iOY}�O��Xբ��U'��ɳ����2�0����F�<%��1�����Y۬y	�#&s-�ຓ0Ћ��}6��t��9�1�������C�W�6n�"y냱Z�qۤg#H�  Ɯ����Yn���`�2+��� S��3�bj.��d�B���f�z��7al��>=���b��(��Pu��"M�o�	�μa��RTq��*o�vOG��妍���"��NM,�?��ۯ�EׯJ�6@����
`3a�`{#���ް�l�| ��ڳޛ�u!*�ʣ'�h�p��1ٲ��A8��]X9v�4.놧�j@�Y�΅�Fο���Wu����]	�6���X���VS�T(��ܧ�����Y�N���m�C�~L�߂�%�%Zo��H����H��L�dX�ķ8K���}7�n�C���\�k^�]�y�mр�>|�X��(&+�H�� �P~���|k6�׋����
�>�ᬄ�م.����>[�:]0�4n.d��k���F=���%�����	�X0�!N��8|-*��nY"�Lfe�/T��٦�!թ	�'�&g~!���}�J��8ݎg!�o� =���`J6涖�.�1�C��eC/�(gi�|�Ri����z�ꉻ��o����d�+|���o�	"6�L��(�̻����J[���^\��"��wo"�
O�R���˧x���``�i�bY�Џ��r�^x{��
H��[ȃH����	xC�k�e��v-�r@2��t�|�M�~�����i���q��on��t�oY�,��~�睅�8���H���L ��?Ru�@Ner����6��2V��#�&t�� ��j�B�O�С��"�)2�˧�5�e�B�ʳ(l��ͯdc���,�����;v���o�,��k/��6y��B��0}���~`9%��In?h"fU�@f&:�2���L�4�z�������h��&�%<�����\����*�!`T�Ȩ��	YD��#xL�B��yc��gv焴"��+h��zr�V���`����
�[u.���l��+�
?w�̷�̫Vb�
Jq
��MK����ծI������F�O�iH (�MH`���r3L�:wS:S~f �jC7^����A� {��q��PJ�f�����|ł���;�a��w�c��a�� ��J��R��[	��W�(�F���6��.{.��F����n>Xh�M˥�)�C�1�f�� rVrr �[B�AM[\XN���R� 1	��i�oy}7���Y��Nt;Gx�I�õ��m�����g�>�lh���� 6TI���ۍ�Ehu�7D0�����;��"v*����B"��)�5������	&��+,���{9q/I3�����އ�/��V`��6a��@r5_O˭��I}�{�n�^�@�_�<�Zxj�R��N�������(���}�]�<6Qu}�~�����c�D=�Ѐ�8{]�l،�/"���X��z�P2����h	Ovv0	�q;L�ݥ;W�F)9s������]?�{���&��^+�2.'+����¢ʁ��-oz�})Q�WJ����׬��/�F��2e�4&V�FO�f��'M7%\0�d��ؔ�ed�6�誂�cOS�a<���]9�XJ�T�x^*/ ��d/�
����t�b��ls���6�g6i�;��"�y'��Յ�=^�$�fp����v����ۧ�`�L)��hbd@���ꮔ�E�5�e�j/q.�V��Pd@���a��8�mr%UTWl��$�D��������F�]X�x
�R&$��z�X�����$Dૼ@ �~6x(߹���c�(���f5ɻQVm��!�(T���"zc]o,��������&R��b�zϲ�U��D��Y��Z��К~�ng�FS�S�����+���(���&��F��8�%:��q�K�.ho�V�������\	�O:�����6�x��Z"�+((�KӀ�J��h��Ou��>�<r�"j��=khcʣK��S.(�FG��������+��n�۰�8��zԵ	�]�y�����Znn��j��-�[.�jw�F�eN}(������WυwD;,��g͉�+s��5�H[�#���WB����!1�{��/#:�L�9��c���i���fz���n%s��o$�������m��=��.%腣n�S���-�ߕ���>���@/l��]�j�<l����;x?%V���$m�z��]m�)խ6yPtD�S{���{��&�9�1M����t�G`�,Y�1%��؋/S�Y(jJx��[|.I��_c*��w#C�� ��b\jʶm�[��`I�N�������N3�����h��Ѱ>�);9}�2xכ�[�n��L���T��������m�pJ�Q��4>t�����iW�u���Zp����e�O�>o	��;����>�*�I�'c��tf�{�>��H�����n�|��w��������/^����^Y�.�	[+q���41uV���(c6ЯVJ>�u�\��8\6m�Y}#���۲�F��%�֭�����"��5�[5� 81.~0��t*]}��낞K�J�dk���$*�8�;<{8H��KDҗ&�i�N�n�q��Q;n����q���gQ�aF>����i��$�<��ކ��l�./��N�;]��~e�:��Ʊy�����𳌇	^�y�_��4�I5V���u����8�=�T�mQ�U=gN=CY�\F��&H+&Z�%[��YSq�zd���/t�����ꗹ�0�O�����k�~�.�;oE�٣,`�p�C����}ʞ�!��4/Mt�4!�[j�&j����CC�?G�
~���Qd�e�z�))�<",.���C�1�-@=���#�����Y��*�"�H�c ��ܶm(ى��0@��"�T؅6�0¬����:$�y��q��>��,ا-q��ˮH��f����z8qdC;]ch����!i�Q��@�qg�YCBB���f�̧�A��#�s��u{��@8m��z�#�&(p7�|�t�]����� K���=��H+hÌ�!M��2,�x����g����I���2ܶw�OP??���>��U'�c��f��Ð ~b^��Ky6
?�P�y���)�{�,�UkƤ� e� ��5��.�|��+zj�MY�hw��|������,�z��Q�!����s4������W��.(�]���KS�˟�7�v_�f��o2�f�T����%ϻ�Axo-�$��.Ι�n�-s�"�/M�e;L��ͦ���+A��L�ժBDAT{U���`
RK�:�����P{^E���7ڥ��(}Y>`դ��^�'W����Z�e�`��r�������ǵ��A��6�&��`������H��!J檞S�z�&vL��^9�&w��J��؛���)�FOO�,����ƥ%+�eJ�����g��Oc�q��;|C���|�2N��o,e-��3<�܆�����#���:�����r��J����B����T0���O�u|�
a�\�|vM]����x��˶�]1�'V�%(��Y*A��ʕ���n�%b���v�^}�9�ZY�Z�����?�#;�W2�G�@#5`�`�4'�/[a�O�Թs�w�Ǐq��W�h��#���$7��7�j��	�} 5���VO6��N9�`�m���N���32����vl���˗|Td.;w�����^��<읱�r��:���OXT-V���--߾]u�}�8�}?E���
�y痧��~��-�?,�D��C�`�=x35R-� ɇ�ŚJ�Bl1/%녇��x��ִ�����U�/����o�y���"'��^8���?�����f4��<7�~8v�3L8��r��.S�~[QJi�{��K�ю~θ���s��0��~�0h��B*J�*2�p������.Qڇ�o�a��z�:!**2�o�����Ń�ū�2/���.�߂?�=�2U�2qc����n����DU��-��ƤܥpR��*�n^1A����Oo�j9���W�^{m�n`iްM������s
K����G7��*�4ͽ9���K" Tg�|	ʑ�6YY�˱�[�;���h���Q�9�k<@����d�u��҄5n%���ƻ(��mch���h�p`�9�����Q9�LA[q�e(���O�epO2A��0!n�f��8~p����[��P� � �A��)(�>��o������=N2��"�/���Ԥ�ƅu��M�́O%Gy�ρ�5__��<Vd�溷��>\ER׷)�J3ٝ�Ln�m� /+�/N��#��A�qV�R�%$߇]$GJ�7Cl���<���h��<��B��
��{��u½|�g�j������u�w��X�1��_�F!x}��[�z�����K̞�: �y�" �A��ƚ��@v�JV�w��+',� Y �yfD�!@@����-/���l�
v�F��<���VnJ�r�({��B���C3���Q��o#A���J���������X��엡ܦ̓�䚹9�Pu��i��˗A�tt�ݗ��C��1�:J=[���ш��Q"���:���N��E�$��6�j�xe�����2��Q��>J��	��/���7͇�q����@i����O"+����oHQA�#�����7��/��U.1(YJp(V�l��]��G��!b���3Z��W�a�:��	�C��.
����_��������guu5$�P�֥����qL0f7��8ߵZ)(���O�̳���P+���vx��ƕm�x�L%M����fR��&��D�xȡ\y>���KzO). �Y�z���N�z��ϟ@Q+3�A�B��\t4�V��n�r��'f#���]~B�~DP�A�8����!�K;E. �h�u��&�Ck�����[%7�j�ع?c�Ƙ���zf�3�x>A�g�V-Ŕ s �o���\/�)�p����?��Ck�z���=��̒���ȓ=��OIC���f\�7?ko׋-�U̏e�|o��U�tm欤, dv��;�D��c:hL����	L�;�B֓�C��1�L���%m~�ing'ũv�!�˿���@v|�e���Ok�u!��9z��xez��h�JxD0�Mz�.�u�wƱ�ޡ¼۴V�,���p{N3�􃠒ݻ\{{8{�r�Նz��eo��8�;��e�Z����[�2o_���Lq�\m���"��U-4�I�ݞ`j�S�8����m�����is�֜��g=n����S���7y����m�G�2��&���ՙ"�K��)���?�n@�W���ya�7��B+ֻ�KWG'{��� .���DA_���[����O4�< $���2O��#���-Ŵ���J�k#zR\S�r������O�78�Q�)��	� i6�(�2�`J<���Vn\���=2�8��7Q�#cc�a��"1����{Z��,�Î%�H-��T�j�#������|VN�s�����=�w��ۅ��֌�LԽB_8��NvL��<��+��;�!�;'��]Lj��}�,� ���a��R�R0Hy�}��maX+7�r�[h+�,rw���Q��{��nY�.0ԁ��|LNQ+�N�c�׬�.��i{{;�EPq�A���W��CqO��������{t�8��˱��kv!��P�hZ{�g0�kB�*�&oNu�y��� _�.�Ր7���SX�����Լd���_��r�HuR+돷d��	>�2�ڡ����57Q��$�<F�@&7o!4C&SM�Ug�����f�.�Ⳍ�P�ڊF����7��CFq���9���e���9qD}Kx{i���[�{�\�C��"����~W$�Kʷ򅷓!���\���*6['#��}���;lZ�ӨSJP��N����X�y^�&+�QɈ�f��@�^\�"*�7�q<����wl�B^����Ug\�: {�ŀ�{(8�L-bv�:�"*'�����LE=����2'Yށ<U*�:8سs&�	���/��S�0u��鑎�N�4��;��+˯�q<8���R�T�mڀ����R��e�J�C�>5�D/��;���:e����hy��0{�:գ��Pٻ���]� ���p��5wsC���]cR`'��`_�l�����;����;�ĝ������L:Ȇ��G{e��j�_���9�d�^TP4�<��r�I��aC.:���u�6�l�g�W�K*t�RT���v#M��1c�h)�<�p�d��k����0��R����'�,&�!Vc��F��a�\��&�Sa4Lk�]6⎅]��|�47I��:��i��UPל�y�w����];d���4��L�8���Cc����D�Au�ڧv��/R�&�X�J붞�l�L�t�P����%XB�l���(������+)�uJ��D5�bf���SB��K7�ߺ�n�7������ݿ;�Y裭�JroW�Ā�Aŉ�&������KWg�ȆU7��'�*n!��:<ِ��yG�㬴��N����7���S8r"g��*��M-LtB����WPJb���OZ[�����Fљ �ߵ ���|���w�R�}<�~t�
�8C���4�=q�h�pP-5u6 ���[��ؼ�E�[�PPV'�bH0�Q��R�=mȱ���3P��D1-p��� �ݟ�r�WW�����%K�v+�X�z�:10�6<� ����$J�*��8�ʆc&�ݔ�#��1hX
���"�Tr0�y�a�6��f��r&a��� f|��`c��VE�X!�۴n9�95eo��_����$� HCb�?�sB��Q�.N<��;%�dw���d9���o�1�nNY-�i�w轢�o�A�OE��=����F��k]�r��<����� ��N��q�.=�u��l��YB�ؗuho;�~eks�*�F�J��2q4 U�5'G�&���N���b%�3{Z�~�r������4~DE�-yX��������- {dd��hz{�D!0�w�l��L�q���~'_�_YA�Ǿy����'�U��Ӛ�/:&6�vȏX礆�'�.�'KWMPL�g� ��'�J�F���e}����㊡�څ~������3 ���x�n��Zr��Lo��OY�@��Xz̷6��4�$�] �&��
@��+��&��Ç��e�l����7��gfϞp+��Rl�dl.��R�I�wZ|��������31(�ʋ�;���5�"_�D.i��w���#
� ����f�����]�I��_P��:��xnC�o��?�Ր��rAy�"�W���ݧw���W��|��!" ��%"֕*�m��L���W�7b� �)��ĺ����.���- a�蜑j��n�zDn&_,E�3_��l�v�tu�Z�,*|��s���@�5k�C5�]/A��(�U:~QT5��9�)����㰌|Z�60Z�%JȠqWN|��T@�? Z�;�8{��K�577����UjQK��U���/J����t@I�UN��V�%qz���)�� ��(8Y���F��..y���<� �ğWe�׃<.�(�M�%' Dv+$�p&j�����r�5�MZ|"�(:dȝ~�e�/rl#��H	�����0�+�f���&���.��CՊ�5�Vko�Cc�+3�Hy)�{��P}]��h�R�b�j��.���/\#��I�>��j�bd������#��@^',K������㦓qg�l���_�Fڃ�O�F� �����luT��O4X(�es���b�Rz�K꺛;lӨ�E�"���|ʸ��(�#V|����[=v���Z�-��۴Jx����E~K���e8�\�{;�g]��c���Xeݠ:i��_�	7Y���D��:�H"�d5${v����[=��xų�m�kЛ��s�m�1_dL�*����f9 ���\�(ˍ<J~f��띜W�ٿ�*�oF���oP����4ǧbګ�����鍊WL�ԸB%��p3�_x8�����q����x�fF��{�8���ݘL�=�Zy6�VRd\��!2�i߫�\7V�ekM�|ƣ!�2�b�^��T��[�tUu�� �TF3��<��{۽�r�]W�?)=Ǿ�wdⳡC��W�k�p��ʃY��e:$�6���[]1��?P�������i��.��X:�} �
�^}tN�O�7��O>fg�'���؂52���4+�b�!S�x��z�/� m�=Կ�d�)�;�' ������$��^�q=�^?�!A֞ȒL�l�ך�ܷv�%ߜ�;�x�/UM��e���̃x(��(w�)�' �6��� M��&��Qm��Ǘ�[��U��Y��Lʞ����'**���v��k`n Z$����T�ou�G������>��g���#ܭ:)r�V)�vS�G���Hާ��)���+�,S3ԫ9�m���^�쾱� �<��wCnl�͏�K:�����BO��y�#r���@ x�G4cҿ��KoU�M�(���@�x����`rt}�ۭٹ��L���c�0��N��R��k�P2�\@$>�hv�4w]�B$�������!��ׄ���&��m &�6Qsj�0N8���<�89M�'L�i�g��1/<x8L��B�/�� �QP�:T��@֫!�q����W�Ѧ��n���5nP��շ�T�e�K���� P��-��3|d�/n�1C�<b���p5B�ox�?��.#�:�7'�O[P�{�K�!�F�s����d�0X�4�4n�F�����S�Es��d�Yy� m A�����m #��x2죈:��YkE�l��Y򶟣r�c4�N�j�ơ�0܍(U�b�@�:be=�8 km7~��a����z?ȧp���	L�qBF����k�(� G�fK-��Afhj_�'Yq�LoP �=c� 2����&KS��2�*�{��������M�	0��T��0��Ғ�� �\�46�פ�a�8���|R�a��mb��2Rjr6S
��o�)�_��Ю�TtH�������-�mp=�ybH�\ ��7�+UAa�`@���n���	�i�w�F�Ͱ�O8�����[��h葻���E�^_$�����ט��^: �rJ�Y�SG����rN|��R�C����w� �j3[4i�IU��ܞB�GDh��E["��V�|�_Je�A�Xt�%�͚u���9
�|_��`�Q��&j���-�NfI����'����^��$��@��w=�K֍��S��_�,��3�6���u|��a{�'�}�u��ѻ�e�̉<b�1C(b��s�m6>2[�Vil�_M��9��	<\*Cy��gUP�d��@�Z��^|yni:��j7'�i`��|R̷ɋ�\�@	$��Ʀ���X�o�K
�Lej����OS��1��y�X�E#,>��y���Zh��O[[[�|t�ʖ�zĩ�o�;��7���ʔ��zES�?j���#���z��}��\F�]��L��FY*/�G����� ڂj�$==���SP:G�G�������ny��7R�K����M��W��V� ����N����C:yS�<wG$_�Z)Tn������"������Mn5Q̗F���wl�"5�����(�^kd�����70B��qZ�ܲ�a�T4�)���2:��rj$�KB��>��/
ܡ��4u��F՛����/o���go�O�9 �T>��A����i��U�8Sp��0��iW�;��_��y��~8|�A5�l��8	��'�)���s��Nj�ڍ���|�SF�s�Mޥ��'���<n0[��N­����!�uZ����1���(�e��c��+�(|R����J[�������yൈ�J/�8;��ZZ���m��p�68hG��3u��@��0�	�E2$[�I&�׉�g�q�4(3j;���Y@ПVW��=�
�h`&�B��
����D��l?�]X���G��{��
��T�*Z�=�d����WN����e�t������rQ�|~r"1�Loy4��Dz�4�Ɵ�{��_I~T9�/:�疝0+Ss��`g�Ǐ�q�݂�a�@�U�@��?�JCí�x���1��r\Z�za�Z(��E�����L����%�̠�Fض-9Cv��փ�_)�oLZY6t�2\yd��1T��F���XH$�.��k}�c����[ԮK}<���ԤYuS�;��-�9�
�#��m��j�;p�۴�R�&q!m�Q���<
S[��*N�ӊAx�Li~�-�*�{��O^��~�\�Fa��O�&��� �a� ;t�CU7��5w��91{t�fB\B�K۔5/��1)p�����w{�6�����Jg`��^iud���Fݶ��R��3}hJ�%AOl@�介�S�ܜ�����Ef��7�L����J�B�P.e��Õ^ �;P���B�CIm���se��Z72��!������"�'Y�6�[`��rs}m��V�n`/���"v���]�U��Y��xm��(�h\4}::S�>j����9�Id��(���i(Ń`:00 ��
�W�/�_����'��{S���y�Ά��{̔�����qބ�����`�r��>D�q���e%29h��^�a�:�q3j����ԯ�V�xv����+�����P��e~(���:�b��˦ nɆn���������b��뺷�ˤ�$�j}}s��DS�
�+�f�}��q��p���c#��\r^��viD����S�����&��A��T4;�Cm���A}�x�����߰딨�F6Lb1_���y�}DͶ-�GK�¶I K���v�"0�@�G�PBSE���T.�	n��.mRt-$G �j䩟U�ޑs��������7�9ܭx�<Z��m��A�^Sw�_,s��'�-��F�i��@e�m[�Fx䱟�L�g�s��s�<���r� ���B�q?���w���M�6��#��/h����� �`G�N��=54y��������M��Aզ���g|�z�c����%Wd�I��3�h` P=ؔ!n����_��)TZ���P@���v���,Lt\�<.��w�����f�
+׹aq�|���z����[:b�3��R����F�9��)���Q��őZ�A�;� �(,8g�~Ě�CKV�I�yN�p�����^Ya�Ǩ}Fjx{{��f%j�����H��z���A2��&pK��D�+í̋��]���¦&r�k�P9hR" �j�T"W�����֞%鑐�?Ev�.e��s�5�ޅ�ل��-7
c5U0�6�m�ݺvݚU���{u���������9SC�g�	��r�(X������Xxb�t�;A��+�b%�f.���N��q�g��T��<�*��&**)e�<��+P<'��x4�f�N)�������3���@�I=}���m�f�۟_�ȟ��CG�����7�d�uW���-����",�S��G���9��/i l<�GTDD��62���y}�wѶl�!�.kKC��7����
��_���N�Ww[��+z��q��#���'�J���� �Qj)���C�޲RW,B�׎G������^\~�*>Y�*�zo>��u
��-������K�0dＯ��+��W��M7��.�_D?+��z#^FG@�r��r�����9z��nSS�v�S�bRW����g!Pb��L+�).u�6��K�=x�D�7��4n��P�k��=E�����jF�#�ժ��$�=��ސ��#�d��oViT%�]`�xC�RzkU�Ű�l�M�tN)QF"��٢�?�b��e��놮����?�rA�/0���hd�?}d�A ����s�U�$h߆$s�im���sB�c�⩆�S��J<����AHs��kR�㭳���֖'��Go�u�ͻ�C7�|7�<��u��FQQ1AG���	���KU�(8fl������B��*U�![���)[D�����~�f���E�MU�����l/��L�^�G��y��%t�]<����)_���,��0�޵�F�;�Qq�En��::YP\�mc�<y033�lRg�I��Of�`�pO��³_�X��@�����M)�8PI��U��NB��9��Ř8%C��v�yaX�6�f`@���Sn�/��NjpO8�X���X����}a]�=/ܐ����m�����ݫF�ۼR".y|�����o�2(
�Ğ������@�ߛ�1;��^#�D)���%[�EV�漩�K@?�G�vk�dK����{�5�;?��j#�a}�Ő������C1�t)#rssӥd~HI����.��y�:�>�_g���%f���.�v������~#��A�~�-#��pC���x�\�2��� ��yK,�<��*0�W��B�D�w��K*�;�ϻG�>�r-���<	�AQ˙[֯:o��;Ք��W�1��5wAc�5 ���k��kwq��rny&)�4�#�xS�0�)��k"�;�nu�$�
���e�����ζ����g�l�4
\ťL{�M��9������E�/�*���b�cR����[1v�Z����*�|�w�ؘ���>K�����u}_&�*��w�jxxx�ٮ;�/?ž?(ix�n�`w~H��_�����Jd��C7>h|�Q�jr�4G�Aː������Ðf< �|��x�����q�#$�<���b-�@��U{���&�g��'�Q����X������D��;'���4��K
F���R[M��hgx�s��u1�F��,��7�X/z�]�
d˧jP4
Xg�.��𐮨�D��"oι��V/={�Iq lޏ��:���&���/�0}�_ж��� �e�+��-��6\����X$:�s�-z��#����&��L���hV��fo���>R�h�%��Ee[�0�����D��*L�۹�q��:gay\Ո��n&3��S1d��b|彾6~�J`,x�ȅ}]6_v����ʴ������5u_�
.6@ GWI�A*Z���9@Y`�Df���s��1��ͯ���v*l�#�໘H��]jU�;B�V�Ɓ��UMyo�,r��Ï����@6nb��㮱k�Nj
�S�S!>&nY�����{_Pt)�mS�3��o-.��7-�E��k��q�Prr2������u@��$�Ҍ+_��M/���@6��\鳐̇���z�އ�W>�`�Z��7�?�4���YΦ�Z÷�.]�"]3�5�����]�6�6x ��PUx U�W֝�O�<�X��2��f���2.oXS��Q)O~ ���FKk�gec�D���v��9����C�1�c�`�{�ۦ/�D|��+��*kf�B�(� ؒx�<��̘�:��*�W�#?R2	�tx��zɯ�˄�=oo��Ĩ�����4tIv���1ј�C,��X��~{�\�s����1�@���v�����ݟ`^t4Ee��G~�n���ZU��۪f����rt�3)�q�e3@w0@ � �ן����FE]�T6��͜��� �]aQY�Rr��I��7RŻ]x�k�eA�q�<F�zP���!A҇��t�;�t��r�����:�i���l�u?�!��b����ɋ��� r��ҏ�=�0ԗ�O�WuR�^&zE/87��>,�&+��c>~W>"�5@X����=,��~�ر��W�~	620!�.@�M7�O�X�胸ۊ���E�^�WOpe��<	>'>u�<T5�5me�'%�K:<��2�����H�&dÕ�<�/Ͻwp:ɧ���~�B� t�BQ�U)��~�RO������1!##�����x�m���&�$�yP�ytE��W�#�}$��~�Э}O` b�B��h�5�ҩ�`����*����G����O���o�T�AH�DM��¯�� GӅ�;��i�����_��4�L�@��?����{���0�����H陪LJ������m^$m����(�(�������Ϡ�_	
v��ߏ�||4�2�i7�#�*�T���#eZ�ݗBg[4+��~E�u���?�;M��`��m5v�Qɟc�6`u��m�ԉNt���:į��t��]e+z�)t�i� *�1�3 �s1s�j��09�&�B����0XP@Q)��=��N��%u���w�g� 	j���w�n'�;�X%�ߎU#��������K���f��mn��t��ټs��v��J%�I� �y�$\���[�uc�b,��5[��4�2���t�/���~�Qq�f�y��ɖsF20BFa�'j�
J���iMew�%��6�w�զ�\K�1=��/[�Z�K9d=$�Sq�k� �bc��. �D��.�l�މ콹���˻ޭ	R�5�������{�3�:LR8yO%R�Vz��r����g	�	�#Wa�rk�^�ZH�W;Rs�`�~b�`n��	�[۵�
2��uF;�X��V��;���E�Ʊ�nǑ��|7����Kn4�0qx�2�
3�һl*H��8p"��#T�L��\[G�Є2��^�3Sz�hhz4}�s��8�!��!��=ExNЪi�dG�K�r=����1 7Nv����H@��uu��� ڍT�!&���ݏ/�za�T�q����u�&���9���x��CR���r ��ҥn��][С�|0��b�&�n�Owv��Kъ<i�
��C�lV4�_��nY��u�p~�10��v�L�P�Щ���q��n!�?D�@8��1�R�N���Ӱ�����P�@޷�����M9��]T2t���]Q�o��'z��,e��$x�6"���ͼ����K�{R���^��c 5�6��W����A�������M]�j�[�-7�W7N��F�j�Dj�{^�J��s��f�䬭KV��6��\v�ҥ.2D�	�Ni;>m#�L?I�9��nyOCHtPKu7)_��J_��9qFS�fF� DPċo[���v�)��9�N*�ZTWQQ����c��t�%�,��?�K*��v�%>�]-�E��{�s�L�l���w�0{۞���k��u�w)�˜�Ka�/37�8n�����_Ż  �{������^ߊG��եP��Y��Y�}nV�	��˽{�{���5��3��/�S\y1�����b�N�0E�2%���ۏ` y#��PT곑���HIA�4ȗu_�${�yy/� t�m�ked��I������jr�o:�JYY�'N�9Ȇ`�/B�>#��ư��p%|�x��Q��qYf[��p�����R*�*H�c�"!! ���� ݠ�`Q�H����t)!"% �t>R�����~���}��Z׺�����w{��ğb�/!3(�4L�J�rq@��Ò�,��YN�/��8��~P��+*��R�S���>������#���C;��ɂ+Fp��YN�b�@�U����.�]��0���f�$d��C��i||y��Z��`+ *�W �og`\u���}=_F������y3u����^����f�v��ϼ�V��Q�ٹ_=d#r��|d�BO/	��Z����$�' ��}�\���mJ\�A���&5U���9A��D���)*)]?�3ښ����tt�Ed	g �	�<
�B�ɦ釩�zƿ��6e`�Zp�á4���.�i|o���r�#]tf���uDx�F��8�\d���,L�P�Y�eA�ys�~��Ă�!^<�����է��n2n%���g��y��(��q�������k#���F!�i���a
����I~���*�U�.R>^��D?)� d��o�GK��aѹ�?+��dd���}���١i־Z�il�X��q�Nq\��'�"�j�����d�Za����I!�N���!���|����cB4VWm����Y;ͅh#�Ј+!��y��`~�Ҝ;u��C�օ�n2v��`�c �I	G��*[���c�?>]������~w�r쏍�8?�9P|��l_7�caL���.e��o1��hEj'0�$%���?N�/Q�W�A���2�
�
�:ζ��^�&(s�MʾfǬ�Q��]k�lԳ$vxK��9=SZ���Ņvj�q�#A �����db?����l�%��^U���&f%��+��x�a)��+n�cw����jq��f�9���ȱ8aINi� �:���=�������Ǐ�4�2vX��>���m�(���R����F�T��|pآ�c��<�\�3�5�<�M<��yR�M��|n���~_�����ʺ��%y@�ǫt�`e�T��k-���( GL
JB�&�ivL~�	:�k�vK�k.�^^�13�t�-e����Vd�^�.B�����4`"<�]��)���!(x��) ,5y*NB�9R���!��e͉�[L]��|��y�ӑ���滪$Wڠ�x�%��{��Hy��?-��V����u�Gz���_L����WڟO,NV�ʘ�౐J�sC�>x�ZPJ�hct9��fmm��f�� =�Ԡi�]�o-"�r��R����ț�'=�����VS��(i�H�E��[:L�����_��@�;L�c"�t2@��Б�����_�_`U�wv����ؔ��J�����<W%(h�U��]�����H̛_Y���$ux�ή�������/mY�ب��p�f������>=>HpJ�q(6��H�(�Xk7�V5f��l�P�Ԋ9`!�CBC�(i���̆��+O��f�h-��v1���]�9`ЛfW��L�#�\S�Y��]r��!��fO��d�;��|b�u�l�UEGGwg��WTq�A���hg9福���6��=_r��5<
�&>�9l����S.��g��D$�T�E.t�t����p\!���hcŢ,xO�R�b����܉@���Ts3��7Р
��V�M�#���Ę٘f��&K��^�4�k��۷��3Z�;"��즳�gk����m���ϕ��8�ɢ�4�b�����0��?��qX���uKk�9��!�Q1C\&J�`� �ņ9�ք����ރ���{� @��p�Q>�F��GHw�Y+
,������/4QSX�k?arD҈[��qa�='��G/��5����HT�O���y�\�\��p�` RJSEq"��Ȥ<j$5�|��"�{��o���wwR4�N�P(/���prFdoYr��$g�y����α��a1�`�G����j-D�)r�[���sK�T�����LWs����z��4@+��mK/���Z��k[���F��@S���H[��dd��������s�/��ݝ����,>ZX|=���̯�2O%H�CNW��*(�AHb���0�����F�Q:��2B
0%e%O��q����I�݊aFFF���+�ǣh� ��ўc�封E�����i+ݨ�ݱx¶��yp0���篸�j#�Q�Q{s�rᜆ	M/�'�.:^}�l���ʶ,�cslsBn�(�:�-�2U�L��K�ؒ2?��������8�m p�������.�꩝�����M����\�4�;6	kn99�!y�M"��S�\W��*�@@�9�o�///���{��D�`��DV��� �
��~�r,j�Z>>��m#ZePvD���,)��/����3t���0�E]$��;A)f;��K���fJRCva*�I�����|@̑����w9@l�v�{�,�^�=�88�K�en�ΰ|F���'�@�"ɲ��%�Q��7?�����Nေ�ѻ`��og|�N^bۯ~5���He��>lt��oNnk��V�m�=�\����R��@�'W�����UHт�r�|����}��]��옃K?�޿	���H���L��?�;EH5ygD�j���f`^��r�����I� ��uʯ��؏瑴r��,*e��I�l�a�6�nл�+v��46+&]��1@>q��Jڍ��v ;H.����Oԓ�6��I���~u�F��h���4o��+��il5M�f�u�"K
@4�xWS�a?&G!�X����m5�ZZ�������U���)���[x��m?׀ڍr��Ò���7У��|eh��TD��u�۩�g���L ���)�ݛ��o�iʥ,Q/'Qk�ٽ�E�CfN�N��-!YV�J��9F �t��/�$��ʲ��eJ�~xz�S5,��y��C��yh��ڰ$�dG�������0���j�\�IB�ל��tD{�k��H��UR2�Wh���-B���ùB�9��"6�;�d-s�,Yrs>�"-О��!}?��3�+�/�!H8�f>r.���w�̷��p|� ��v�X�������L�"_���B��;�v$������{�<�2ov�O[�"�����f&��{?�Dه����q��2�ha�4�ITc��N�k�]EoL�/P�A�bd�n�r�q�F��	��#�����l���/\����Of��l�)�� d��ȯ��A%�-y55��u��u�u�;��S�1V:�yO�9)��EeFd>\��Fz�,�b�x%_��<���wfH����|�h��3��0&ܑ7��H��l��`_?/ʷy�Y��Jx���2/cs����,I��9�E*�J�I�E_����� 
ncc���KI���������y`L��^��IW�L���}/by*F��4�l��g��S%����<�g���CJ3O�[Z��5��$h��:LV�Ի�W���|�tX2Һe�늡Cs����c��-yw%��,26E�:�0Ҝ�
��7��;*�	�wOyG=�!� k��OxY�-N�^ݦfP:?|���c[�QՔ�w�i������1B߂`ZmWD�C
#-=���ѯ�֓f�#�4j�Ә�~��&0�2$jd���"<�ԑ�d��I�^t�Z?�\G����q'3�e�*�uk��u��*E;=�N�6��t�����d�JnC
^��Lz�+7ė�����I��<=-e[��CǸ� �R���^ W!�V	feOpc����v̚ۂh\,��%�ڄPOz[��d�yaF�X�����	�zVSy&���ҝ#��gee6o+�-i����`_��ƽ�b���wwfC��������������o$m���X�Հ��ҥ,�Tn��')��I���Tr���&���ÝƲ��cR����hhtk�{���(����~ץ����C�ny{R=[=^=�\8�T	�����n�L]Ĳ0V��ba�Q���2�_ř˟���Ӛ�F�c$�Z�mLm??���DL����of=]E�a�U��09]��0F�Exz��n��ݘ��]�Fܳ�X��[9]�Wְ�����4��pC �YDh>�]_�XN��q3']7�`�옷�d�U���za�����con��Gޡ,p+�b%)���{�|����(5��ח�4S��G���c:?�p3��=���@��I1�y��f�j�?�8�$w7l���}+��}��G"�`M{]�E�cܛ4�
:�L3��L�P�A�q`b)�>.޷�a��Vk:S��\B�(Uܡ�E�DT���م�A����xn���Y�iۮY!���T~�>������	X�x��\͞�*��b{�!�z��!D��u�<} P����Z�;�-�*o#��#\���/k����ܘ�Z�!�X�*�GqY/aʑ'X-�x�.)'���?����Zy��,Xj-�f�L&u�ؑ	,J�F���	ׅ��c���
@4="u����p��x�ߎh���Ǉe��r7�s���ܫ��&��$a���1f����.Ї�UZ����{�ßo!��q[�u�Ѯ<���s���u��=s��
���NW-Q�݃F6�A��r�FF�6<ɪ.���߷۳�����i��VZޝ�p���M�Mm �/��Z%���?AA��}#�Wԛ���H�Y)`d�v�+��ӽ�N`/�p6h���ٔY.����u�b�r����KY�A���Ʋ�P�����.�m!�+}�$�h7��ܨ���9XៀqX}��kcN +�'���z�d��1X!��k���m�<��:PWoc��4�g���N�y����̡��9�k�$]�7���#Uv����m�j\W�^��,�JE`��Q�T�oW��A,���'�|=��'��ChRK�denњ���8� �]`a=�1��:������̗����������k߃�ۏe��a*�'���U�^��9�g?��Q�>aR�b�XYYy�[e;]f�M�w�ߑ~B��r�@��h�����Dc�������0��ɫG�_^&��Pv��ݻ"B��R|�B�F:�o�+q��e��O�\j:g�^��<[^�����/����'C�O���l�/v��Xs���%/�'%v�©� �啾�n��@y⑕ҷ;Nod$�ؒ[��{��Z"�
�X���3M��2>YG1�����#,+aR�ķ��]�P]�˅�����b�]E<Kwv��`�U}�폖�����]�ew�2s��̕i��+}�����A��E$=�P����������M)�Γ���xu�y�D�N�#8��͹�0�@�O;�ߣ_��V���$�A��+����*3혧�쵦�}8�'�W���_��9l���U]N����a�)*(�`����@+�����׍�} �@��M}�ͱ%
��S�����W��.N��4�1YB/��vP�N��[������ޠ+TqG��
f���谰fP�ll�n=^���4n�,/��	X`V
�e�{du�+��NsZ#F�>"gr0 %�&T��T`Ӥ5�|� �/���ϡ��/Q�r��Ή ��7=�Z)�}��.�C$�	��z ����-A����\mz|/z��{�9SZh*����Lڞ�q�iA��S���YH�H�b�!�a�IH#������Tp�09=�	�h@r0�=L]%nNbZL�#w���l�)�S����H޿ؒ��d���m@r�"hw�i�)�̋�2Yo��jk@�{`�������1<�L��l��$H�nT�vM\���y�My�Ie�@H0��Vҭ\�k'H�yOTF�#A�W22�խO���w�e��(9�Rn�@ꌧi���!=$��f"�7�@�!�5�4�8\��ԭ�a��f�f��ee1W�߭��>�܄Fo�q����|�TY�+�*"}d>��Fms��f�Oa��B�����%M�t~�ޭ���8Hkl:EM+
�+JÝq_M���d�-0"�M/�ؔj�[���VCb�h꥿�z)���l.�}��<�G�H޲}?�f;}�+�⥥s�W�y�h--�����ZF�(�~���?�n������Џ,"o?�Jk��,UZ�x��v��茍�U�N�k����s� -�Wօ��.;��Ӓ�J(TO�����n׈j7+Ò��o�;�`��h�5ګ|F��@ui�f"��lي��*����]��>��-��y�Wfq�㛆/�#*E���xN$f��d�����ׅ��
Jj���_gV�5ԕ���
��֕�땪�x��������b��i�)dyG����u���v>�Z��<!�)��_���Kߴ�����^��n;$%*^c�2B/���,=�����8Xq:][1����/��H=���:�|_M�����	r�b�4��"�����	(T�&N8p6&&�gE)\>��6���L�D����]���blC�y����g�A5�4�d���%0�2Z�Ӿ�ʪ(ڀ܁Iե���=�A$�u�5��	�M�}Q�d����NY������B�-���׻����X�j��a���)P��뿇�&)Eˑ�i��an���+�Mx9��tN�M�H'�0���WJ�9���vBt��!����u���6#,��G
�j�\�vm��@LU����r�sq��ߵ�;*�cb~K2�������9mgg7�������ű«�yLxKFW���ƞ�K~G\�dl�g���]\Ssa�3ɿ�ߨ��+p�LX��|�~���(���j�k��-�Y:i/Nz\O2��Х��}�7��V�.�����zX�3�LF-�^9�ir_������2�4�,�f�U�4�ǩ����ScI�i��y@����Q��NHvNN$�Ʀ�Q;��F
��6�b2/�,]}��O)|6�C��>���$"o;[.*�I���Q��4�t�b�q:d�&�PE
�Ν��(�<���2�nrfܾzu_�������	�J&�+G(7B���I l^>�{xG�r���"v�]��&?���v��U��S�J�+�X�^��d�Y��X���ȌQ��7�������[��Yvw�`}}:��,�v|�8R��ق�%[�h��:ٝF�_]�~6;y�١l���i{�N���A��޽
-َQ1�%7�8V80`r�R �nC�ve)_\��K>>��F�:��S�M��
y2���koW}J7$�<m����A^�ʥ��.����=�w��.+�bUC��}�I��f��� �`�8X,��hF&��h�#�������2U9G��YlK)���^�#RR��K�E���	/������1��/����r�7�>�EP��&�R7x@�p���ano/�s�xj�#CYF�t�f�zc�жc�*"�[�B�x	��1E�¶dIH2��Jn;_1]O�<�5W�C�=��G_�
d,{���Sڬ���-��mX�K޴iSI��0�n��{����
�TE�b|���"?��0�����|�	w�g�.�F#V��&�>��l'{�7[�]9m�Y ��%����[�6��Qr����,��2�DZ���\�����_<F=����y��۴�=(b��Vbx�F��[u�����H��\�c�=1�@{>�@_��aJ�'��!U��q8�al�ȑqz��W
s�v) J��9�=��~@Ѩ�~��N�p�v�)6�}T��f|'����`�*:��R25c��>2�&C��*za�`'$�̟�v�Ŭ�����A���.��,,�䣞�3�M|ؠ����	w[�W�}����
�B���a�"���`#�S��Ĭ�ج�;��£���0X�^�HiYq�ۄ�g�e�c�TI��
�4�M�+s�M���8IZϨ�PDr��ў�����K�w��d���Ҽ P�)%�\)���!��/**�^��}$�>/���G��;�l�v�˶SW�6�������D�w?�Ea�r"��u�K���v,e�HD�:E�tݤ���]Y�M��.�R�,�t��'�����n�|����^$e)N�E,�{��8���-_����;?-�4��߮�q�f��%��ڳa�%$Z�Flww���5H.1m��{�r��I�!l��;w���7�;���0L���O��k����9Ӟ��053#���<�)xLBb����:�) �)^��7���{��г���Ff��8&d�%�3݋Ǹ�n���$��I,���k�a�E��(��-X0��=�g�s@��8u.�����n-����z�Ny����� ��޹��G�AR�)e���r`�ᙃ��r�>J$������CO��B���~��Y�|3B�7'��t��1U�����54�pqq��� ���OOPaxA�t�ڳd^ }}�x�6�5�L��� �'&n�F�hfE
�� ����<��H���>5>&��hE���4���Uss����j�'�c̋�.0�ќ����L��B��;��<q�̈́q�d}0&B)��<h�ƍ���@�Ѫ���e��6�! #�w+&|�1J�9ި��/���Y!xF�X&(qp+P�,l������"bV�
I|h�)��ՍQ&A�e�V5�T�X�c-��f�g.�O�����F|�!!��@�xf��4�����Q��7�2��s,{��f�>�pbeeg�:������a������
��NzT���Z���x���@���-��2��}^���]�h󪲅��\�֡�1o�V@�7qq���uј$B1���d~��
~�F��y��#;[��x_|��j�hw��v�+Gl�Ϟ��k'@�� L_�a���.�I��)�l�w#Âa�c�O���8��-7X-�g.�BCp���nX8#{�9� ���HE�ջ�28!zޖF�{::\��+c�������h��ڪgnn�]E=ѹ<��S{�S!~�VLW�7��$�,��s�wtt�����\�c��{h4MVz�\�=s����6p�݇��===_à�����Փ��)���M4'��i%d�t�D�tyQ��d ���Ъ�<7�!�H��*�1D�6!M�d�ک����=@Y�e"|�#{����۱?�5��-���T�R���|��cf~aA�g�祀��y�> K�I��¾>&���#���jl�UE�h17O���vWtt�	3y���C����;x� V�H�G�Gr�����[G��J�op�m;�a�g��ҬR��=;����8��B#�@�c��1�o�n+�+҈u��7�b��8�SH�*k�WN�G�����d�q�����14Wֱ��lM�Vɢ��˄�S�a?�]����>�촶�����*)I�F�6��fؼ�4�hn��N���}�\+QT5��?�:�6��t�Tm�D�F>�v�3$d�m�V�fb��<1-M�gv����]��������JryW�:hh��x�UtG�?A�"���3����p�6��\h >ؒ��y7�j� %�)ioz���6�i��K���+�c��Qe|B!�bء����*����Փ��B�Wh�N����K�������'0ݍ�6��L��?N7m$P@�1&��%�'�FT�(��	:M�?��2���U���}�����k��� ?%����U�ꂉ�����������*TcҰ�R�/J�\��#pB�1U"*v'��T��H;~������-����0����=@}	��
ВA���>����=�F`rF���1�E�|(�SE��m�@����6�C�rtrR3vV
��|��sW�;lX�|�	_Aֈ]�3��i��?b���q!t/��[�����m�xs<�B@o������zu剷�� ��u?�Z�L��[����?E�����"f9f	�����A�8W5���>�jH�޼���y��h��OW����P{^��$�"�:����X�p�`Oqo\����`dQ�Ճ����C��6I-'�bd�-?T�e$���##����Kg�b�iy��چ���|.�!�m �ސ�wF���{DpP��q�%)��V^�́ժo��XҚ���:��.���w,�#A�<� ��9 G҈U
�G���8�0F�{d�i�6��J�0@^<�>�O�LA�# 6�����=�U��r�?��Z�?�`c*\�fFR��v�A%����� ���zК�;6��?.���ۢMS�(3c��%� �*��-F[�)���g�hy�f3��Խ�6}`x��/��:lO����Q/���n�w��bn2|��2�W�1��*�V&�Tَ4�Z&�SB�!x�{��E���b.\�t��r�;�%�N���m�����A�'T,��$hhG�=�y�hܔ�]��������rG�ٌh�_J���^����.���ܙ3�Z|�Fb՟ _>-`<�٘YY+:y�鍓�'_^0�j<h�H�[0{���~?m��7�g��I,ި���������I���n<5��1�����2�.ށ]��_�����
b�,^D�>tE��X�,�8����3�����Zئ�_jeq��4]ᤠ/��C0����2釉�;���V҆�R)�]� ���0)�d`�i?dsO2_������)E)�NI0w�%Q#]'�|�`�	��Yc�j���eה;�3I#���e$��r<���x�&KW)��Y�Wa�+��B	�;<+vF&B9�n��'ɽ���&���{ϕD/�����L()�hG�3;SE�RXx�WY�P��k�g �M���\(/	N�W@�`k�2xz�{�&���=	z{>{�Ī���x3]�DnS�5��4�VQ��R�m@ං،T�����4�`L�&���{���i{��S_��a�W/1�O�]�`o�w��Gц�ڒnj�+�D8HX��'f|�v�'jj��>p�5X�M��� ��|U]�B��K�6rG��b���F�0�#""\Y@�HU�����9�W2�\[��)���1�W�����梩f�ٙ��D��¨����m�)�����
�Qs��+n�זC2���������.?�aw�B�:����L��6,��w������x�VS�O�C���YԺ�=f���[00(�~Orr�2K����L��X��{�K�
���cOR�-����� * �֭�4�t\&�]�� ⛅O�
�ذx�4��f�(�߹uk-D��)���� 8x���͛K�*C$]�ª�u��}qNN�L*ku�\6�fJ�#��=(5����Z~���WBq�����/_qv���d�y4i�RD�Wp�c^�R[�T��U�q���ۏ�F��	Fb��ѣ�\gÊ ~������7.'�~~��3�1Ug� BQ�n�/�i�_`�9�O�I�[q�yR�~���H2tv��/��	�e(.��E�6�!���Pr�L���,���v��s�;]�b��z��0[�G՚��U��z�?=d��-#����\�2)2?�N���ÍIxM��s��son�[��a`�c�ð֧�2/�L�����7zA�Z?l�+H[�vv1U��۳m��W`�'o9v�ϝi1%0�k��F�b��zϟd�qzg�N҅�{aU���LR�`�`���7@��T���M����.��'D<yUR��o>�=�Em��?rL(�L4x~bo���(w�����6r�N���I�NEr�B��8m���<%��[��'��p�Iw�/Y'7P�%�������x�e����f��Sw�и������;��Mu����X����Ζ^�l���t�ȕ�����3ݎ����,��R��^GȪ��n݊�/`104�_��k2�Kx���8�n$%)|�Þ*���m-�"�zX�R����.�	�Ô�2��u]����v=!�`0������ß�c�l��,K��i����"�+��vc�I��\�4P�:3SϨ�ÞH�L,������"r:J�8_�Wd"tfEF>�L����� ����p�����$Yq����$V
�C���2 XՄ�)�t?)1���B�B�b��l?qq�7��V�>w1���n3O7�W��@x� 嶤-Ex�*��\������[&��7� xE�8D��G,�h~ZNP��M�SB����Y������� jO�QbN�e-���H������ `%��`��8��d�3$!����}*A��;@�G�l%\�.؄k�􉲜�<^?W(~�
�m.��<[�	��i|a�.S6nKӤ^�T!KכvڢQ��YM��a�y��/���$���������6r�b6�7f�Bv�'��í|����v��A�h�e��š��4֍nÌQ���K��G��,�Pc� ���ާ�Aߪ�����`>��q��"�Y�� $�ԩSy��||"�rHp��vb�@`�1-�����|����ĭݟ �xR;��c����^����;X]�����%��D��
�MF$mdl��~B�L>��&����&��0H�a�)<
���O�W��׫�5��*t�=? @��yk�E_���욨�+�q�uu~i/!��&�}K�`��m��ok���iʴ0*�΅����{�f��07��J��w7[�t�C?����,lYdAp�s��I�ֹM�F	�
,|����=������6���.�2���5y]�֮X��Tj&�d���*��:,�ȏ�9<����%u�.j�]�v�e����a�g��5m�N������jٖb��_�� ���:�2�=��@\"���g���KՔ��%��|}�fh�?FÂH��'\#'P��4IF��?Q��ٵK���<��)t��SXTTt��<��6[������2��a������ק�] SB����a��A.)z�9�p���Czk��X5���R�:����Ae�]���7p���
g��a^���C�����7�?�J���_��K]�W��G$��t�6ƪ��C���槭xpU�4�ʻ_g��ϱ./u�Hs�w�{M�����ux Q+��Ex
�2)�u	H8� S�
�t�/�7(_�����SkQ&8�Ç�Y�\+K�Sj��d9~u��\�q��VG�8ѕ��sr��ج����֔��\kJ B��
%�ӌħ��u��[�-MF>%v�y��^�ڗ�<?�4Bb�c�����aEz�Ios�t<:4-7�_lҮ����!��Mf�?��_;<Jp��R����x�w5��/��{� h0 �AJܙ�C�H�%����"�y��$� "�òt��FO�q����� �:��(�����<����]�W��>��.�LSK�,�|�o�����9�M� ��<��*g�N6Z��.���	����ծ�|�f�/�{�t�X��?��6»���Z�.�w���tϮ�.��Uu�����66�%� �Dn5�3��tU{�g�T�{2�D�E�2y��؅m��MN?u�����Q�U��<���c1{-�]]�!��t�zuz�U�<�5V�������R3NLL$M�"i˙!�ś��2K�� 9 v̆�u�r/�zI=H��u1��͕�0�т,���i�������b,�$*W��=�@� �O ���q�ͷ_�
�I�8o�z�VK�!�/М�S33���0�od&ӜMZ�AfھZ�G�lW�5��ķɥ;��V_"�v�͆��z�~ٹf�,�}#����ov�WZ�nd����a�������Ӊ/����������arP���,Tc l�tf����`�r�4ʋ��QO�ż��b���>H�6>->���C@j���,��e�}))�������o�myt��~�$dvq��^KP�L�'�ج�m�W��b�p�O���Y6��NҪ�-5���G��NM'����j�J��J{z���%6��r|�r[����f�����Aڡ�,���f�C|�y�w���/o����޼sl+�L�� *^�n���2��%K��)R#�4���2X6��֏�}9ߤ����+x�2.�abZ�,`@��4T/V���%]c(a��7<a�f�邚ȶ�S�XRK�QG��a(�3�MX�)S�č�:qi�
�����R�v�ik��rt5�*��'��v��aǘ�.�]�/ΑNL�C���:����[ Ɂ�sa������>а�5��0׈�/�*֫��M^|(\?QH�P�`����Ç���R&OA�cͰe�5G܁}�eD�C)�#6�o��`T����l�����y����@�!����x�ei�5��v�lW.����
���	WApG!�i֦v��������L�"���6��Q��ӳ?�-�Gn,22RE P͸�PӲ�eݲdH�K*"���c�����C�E�v ݸ; ��]�[��?�~�R���nA��OҴ� �q?"�thy�s�dn���E	iF�hrrz�2KM0:�@KeW�3���3LȚƋ����?.V�Bp�x�315WE���3r�\��c�/z�~>`F��ggٽ0��[��N`���S��P��ʂh��>��?ءw�(Z��h0���)Y�399�{^hrE�������%��"�������ץ����٬gGy����j���]Җ%&�	K��MCq�ef?F�c��_�빟<�4�����o�0!k��վ�2�7��2�s��`��?^�J5Vx��J�c��Y��lI ����	=�@��e��!���o>*C�<r��?�h�-Ja>r7ֱr��������S��vE�m�h��9w�)�{��]��_ʿ��߶la.׬��#�UbXG<_���d7�h[��y��7����$�rcQ�3���J�q�d��:8k��n�Fe�� o>Q1�HTR����z��ʪTzeeէ�Ƙ�߀_����b3H"�yg<	�N�%i�Ƶ����A
��lŚ�z�"ۑn��{����~��Ƃ�*1L�򆽎�h��YDx`��Y�^ܴy��#X����w�B����ğ��mt�R~�r�����+��y\����j-�#��oE�q�yze<�q�&��DJu�Ԙ��� &y�R�,f1x�4"��s���29vb-2u�ϗ�kע�'9�v�vt�]���G#v����4����	�;+�Ԟ"�_x��={��H�c�^��Xﾚ�D�ۀsC����>BySS�=5|7��Q7�R�����i@�'+ӳ.�g�-�BWE�ZѲ~�,�9�ng���=:\�2�;!3$k'ç��ꂠ9�Ֆ�硝�툛~~H��kݧr3f�u�8���^���jO�{-��o��v���@V���C�&d7���m�]����ɑ��Wó/����qi����W��d�nza>B+�e9��lm�bz@�;��o/*\����RO{� �*���"�y;�HY��t�I�mq��T"�K��t�,�:Zl�dd\�ZZ�@�:���콵��$t$X�_Cҫv[�$͝��@@��"���U��`������odM^(n�V|hx�j3�@E
���Z�IiF��U?l�{m�j<����+�~0s>&���q�R�yk����P'D����Wc��7~��⪅`I��ɧ�6��'NDG`��>���%NNe�8$`�x�$˗��� �Ng�ö���px�4GG�վh󪘪{�a�xyy9:���t�����^��O��_B] ��7��#|��B��˿�W���2-�����i�31�0s����T��(��u/p�`	3�G�[�Ҙ]����`/��o	:���	��Ǉ����rz=�N��N`n�P����j��x��\��ҵ{u�W\��މ/����v��� ITh���C��� �1[Y��)|xϞ����p?�J��d�G�n��&��mYV���7�8�B��l��4���T;0�����~�ؚ�Tx3lV(u�?4!����f����V����
?�=@���;u��e��ؑR���yٌ�kƶʍ9m8_a1�A�ѳ����s�� �Y���9ݤ��6�f�T�d������a1����Ax_�����^�i/ͻ��s��3���@`
f]�Y^���q3������s�~f�����8���ǹ^:��_k֮7is��sj�)�|�mq���Mw������ռ�}Z�@<1.��fz����i���^D�����R���rN�Ä<�[�M8��f@��_���d�� ��t��ޮ(�����_���_#R�O[?mgcS200�_p4�ʺ���m-)`���D����0̰3���i�F$�uUXn4pk�$3'}�	w�}���bڬ��rcmO�'{ܖ\��Fg� 5�X�P��?�l9�FUj�Ȟ1;=M*�Q��$:j�QUA����x,�mH�~�+ى���сr{'@%	*���	�zp X-@�8����C�nq���#Z�����C�R~�L:
��:W�ֱ5�����c�3�?��^A�1�v�x:��x�E�r���	F5��X�.�����8��'ؓ#F�qc+�'�" *� ��T��~�V�<f-'�:�7(]Y6qsv�Gs�N.ߠFq�`ǆ�y�6_	��c��9]�D�ښ��{�Z4��Ar\1����M��ã�6~��l]���uia��l4т����9�]v��=�ѕ�7�k�A��JQtJ���|ie�����l��ů�ܾP���D=^�D���,]o�dQ����)+��řV�?��[p�hZ���o���Kc�Q�@�}��Y��P�����FU
��h�2���xg.ʄ�p�R�� ���gNoA���+�����g[J��4rB?���X�Nf����Q��7vyɱ���,-����-�q���e��:������xX%q�;:XCfaayT��+x[zYĲ_��J���,c�t���1��]�(W��} ꖜ�Y60`�V�ø�:"�T��Q_H�o�N@�����iǡP�hX���X�Uk�AG�<���V\iC��+�kp���)+�z@ب���e�X�^yNN�!����[�WZ� �)s�ssW�e<W��&���,l �ucc�t��-ȭt�����U �.�g]w��e�Z%�G�l�IN"W{w���jQ�xL6*���P�|w��y,�~�L��Az���zÇ�lj'\��;v��m0&�%&&1
.�t0v�ZRE�]�䴶��6Ņ]llؒ��׀W��p�[a�=�l�y�Ȯ��X�|8}��@^�*�z��ږ��
sW�9a��̉I�����1!��%i���� �ϰ��1�4ܯ�V�h�����8��ݕ��Z�\$i�����a���缼pزߠ�<p�N��g��<pK��{��s���x����E[g3o�Azz�pS�
ox��\��[��Z���}5�w)�&���=���9������ޫ	x_�^�>Ӹ\��$��߻A؝�j�����k�I�Z�mڷp������]㛛{�������ݗ����;�R��~^���/����&�e��z��Go����(�Cڕ���4�d���+�m"�����B�Q��c^|���J��׻���BB�`�����ɰ񁮢�\��A�/�;v�<�å�������sp'{��%i�����tZt4������?8�Pe���>lQ��l�樯�M����&�?��'L�g��Nxz$��fUد��z�Å�A�q��ә]
 _i;��ׂb��r�&/O����g���K����9U[�j,8���Y?6�ћ���H�E�]s��=x��eJ�ȧjr�-AF��i��˯�s3Z��߹�ٿU��9��)w	a�-Z��ˉS֔�i��y��x���V�wG��G���b&=n���j*o�tPTT�Z���J�w<G�w�aL��s=�A����}�Z�2d����ǞkE�d�W}���_�ҡX�	E����t~�K����#���*akN^ay ��i��O՟����q���w�|�n�ڷ�3&?�p��3L�M?O_pD��ʥ�nJ&H�b�9J�ܥ;��'$�Zw<�}������c�~��s����Lѝ~o�����=���c;85X��Ln��d�o�a5�G̛�q`��`\�������ԥ84sڿ]>���汗Ns�]ͻL�U�/)Ӑ��1&_Y���}�(���#nǦ�=;�+�X�_�pџ�?��K����O��8���w�w>xI�v����I 5Xܟ�.N덜�b:{U/�o��9ⰵ?���>�{�A���9N=���B
L)�Ռ^3���wa��gnf�5(N��v���-O�s�x�=hI7�rf纏����W?j�0>������/e��-za:�b����{�k��������5ΘG��5ȍ��l�vy�V�7��1&�_���j\'P�����
;S?�m�k�gbb��4pu�{�����8u�FF\#bMk�Ӵ����7H�H���J��@���٤������`���|Ϟr?��̣�����-u���g8�K�D�]A��#v��_Ue���+��y8y�,�k��f��l������o9[2��%EWռ�7d�j���d�CSk��w�9̤�OoR�]���\dpD�C�tD�p	����_�s��I��kM�7lؐ�8�6��z��܇I)�G�v[F�O�2;�����*a����g��fh�!����p�'�r�˧W}�UH��>�rwE��cU���6?����0��qk݃+�Zo5�ut6HV��L�n�������Mo9�x���1��^��?dF��ҽ$ey�I�i~������G�!p����zS��)KO?��*��/c6��� {�y2F)LU$�Ar<7���� ������٤;����8��<=�����w��eFe���[�Ԩ���M߶�%K��(o����7}�?Wi����Y�����3�b��W�W�d��9mC_�UT+1�}*9�奤l���'1���Й���aw��g��x�x+h�5��uKD�nc��$��W+�z���K;N����r��
�g��A���D��-��k�v&q�m�-Uˈ-=�Ƨ泵�,cy����>x�-���~:���yzp:%{����gk	韖N�j+
��=��b#O��*��𒳡N\��w�4j+9"vҸ�=����uG��;"��/�V[['���	�&I����s��ǫ��6���`lM���zIQY�g�3�iv(�?��u��˻�i��.�R@���oUcM\\��9�������C�*:�����a�+��z�Z��G]���(�LO�tsVAd�id��L������)σΪ>���O�ˣ/��>����
�L�����=��e����ۼ�,3;�j� �?{Eo3S�p�F����7v����o�Iφ�-=����/������4ڜj��0�.�6�����R���p��}	z�jit��_��$ ����!Y�������`~P�m<�2c���8�$�k����x�n	Q��޼3YKA�Z� �����\�յ�~����t���<mӮ�<�9���7�x�ݹ�7^j�F����|Pz�9��{�ii�+��T���:��>���r����t�qю��M���A��בg|�s/p��!I�Y�G=~>>��'���&��g���Zh#��\�`LؽyE�VU	��SJ/�r�@k۬7���v���&''S�L�cZ¢������;�ͫ<�*˃�lb/�b"�1
�4�����=�I��= 䊨����,��ߨn�D_������p,����T�$IFG�
��le�gvvFh����l/�+�!!��MIVFF����}_�����s=׹N�����s>�w<F8DM�b���~<s�%��������Č쨳�S_S����"֓ٓD/����<7	��<����Q
m����hC�=�K�~\K� Q��7=e��{:����*-#�iA~���}F���hD~6Z����>��IG�:�������/�����b�2�ѽmQPD$�������@g�@�ӹI� [+Oi��L�� <��L�zg��S)ޫ�G��=��o�����ks��T����Mon�0{s���-���Or��h�X����:������r��N�_�
F�sTA�9^%���f�	�슌���zeBu����������{�K���oԉ�B��=��H�.O1F��`��Vj��~G��T_OQ����/�[(�NVp�b���+�MO�w�/<�Yj��C��Z�����b��ϓ��n�.r�"��"�_�$�IJb[����߅�����Ӑ(\��9�vs��P=����oԅ��F�B�kK�n��L�P]Q����>�}��R7�
JK �x��?=%/��V9p�'�q7z�ɉ D��Wo�{���B�}�6!1�B����)��|���)������mm7��4�Oy���5�T7��`?��8z�<T.^�(�}`>�m�sm�.^�"���_�!��gzĚo`b��־_��Z�������c����Vy�-)kG0�x��,��fa�#��	�iߕwB5~���^�Q��-�8����s��P���S�"��c���5���Nc˗��6���q�}�����pl����9�i�����n�����h�b�2~��'u�Lt���@�h��q��06��Y�H��R�zg&�*����)��1��)���	��o�OIVqfLN�%���v͛�{�g�����i>~���"�{��彩A�נB3��5���k?��sO����f �L�����I�����kP��U���������U� �Ag F��C�k�]���M��������s?�kfr@�:3_L��W�'�q�B���`T�@gg�6ɕ�J���G�D��3I�-^I}}�?�����
��jL�Ŀ|��#ÒjR�i��؜a����z����/7�gU�6��s�,�s*Y��Y�<��:E��W��P���{�����賓�����߬�!p�C$Q�nN�W�j��Y����aGʫ�ˣw����{��FMvq����Xx�E;!G�^A9�p�<�_�mp0�������''�B��|��!R�eN���}u��_	2�Z�p7Qx:1^t������f�&A���,q�ש4ҹta�%����p:����߮��<�
qz����bu퍊�D������Qξ���݇�޼��*��K����#��:$�O~{�ܽ�@��!�ԏ8hC�������{F��L���Ui��k6�rZ�7BЉOc˶|=e]��Cc�6/�D�H��{��s��S�vΏ��~*ė�*�����.����aA ��C|\��Q1|��9K�e
ܙ[�2<-[O������=�BK�����^*,g�;��;�`�����T��cK�<�Q���D1��t'vxH�߯��j6Zhw�`�6�-��P(���K��\?�.�����{�K��4<�Ć�,36�}6�����2'���y����������|q�}�&�ϼ�ӦW��Ry��lB���)�	��p�4I��/�c��g�M.���&k�(�?(N����isy���Ə"Zn!��{���:��Ӹ�����yj�P]`]r��O����$^B��+�A�C�,�iѨ�o�y9�$5L��#�	���zc���_��`�����_�ec��W/��1�`�>����$�`������:�
O^�SG���������f��L_�����f�4��H%v����/����D�|�F��k�89S��N�1��]5��:m��!w~6�_ ���q���2�MW]M9LxAQK���l�0G�J7Y�I�~]=��CJ���p�������Rm�D'YG��q�YT������6'7�!��f�Kh_T��]M��|{�o8����EMI
=�����_����_�4~?�@y�%lowp�c޸��S�F;���=�g���z����m�����w_k�jre �rӆ�̷KX�.�Mod�s�r'�� %ѻNb^���0\Z�.p������en�=AnR�lC<	߶���x��LJKο*!� 1#�U��M�cHW�9q~��qΔ����Զ͡��L�󝕄7U�'2N������Iݺ�"B��(�Hcؐ�cI�}�R\�C���f�{��t���
\�?��ü��;��P_��QL��X�{�ɵ��j�i D��,�[�/d��hO��9(���؟}(Â�?���uʸh����N�r��a�����'�����sE�ox�:�[��5��Kr���i;��;��;�)��w��G��	�~U{��9?�Sx��v-Ƿ*�p�+ �0!�1��묐?������]��ݿ�xl���G�|��bhl���Im��� :,�q���$���_�o�
��4ϝ;�,�9�O�0�JjN</|�^ۄ�\.��:�ȥY�B��h�L{�����1xE\.ؠ��k,c^�������V�7�^o�/���$�{��}�sR?�h��*�����Y�<��\��d�5֗����7S�>�ct������m#��W'P�p�����z���TI�"~$�C��~�3>|t"�6Y=U�nʈ�c�`�h����@j_��,���`\���X� ����c��qζ���'Z���6�A����d�6�o�=˶����&Pz�,Y�⟠�����P���Sh%*ɥ�Kr��[�xب,�J*̚�����������9h������v#�<�%B@�{��鹶	%�?yT4!%E���T�h�V� M�J8�>һs;3��I	י��鱵�t�]���ӿ�%��cup}}��Νݩ��_|�!w�����"sߌ�{����'t�8=�;�a����h@�)bzi��u5���J/yT��C��A��8�!G�Z&�*��<���7�Hdй���i������O�l�����'�ۯ���}�;y�Vi�M�b��fT@Eo�Mz�+�d]�v��d'��<��|�&�����W�v��W�Q�TU�{=W��<��ɦ͚9A"�X >����neg}_�{Z�]�'��e�0�#�^�r�#:>TS�co<(Uy�QP5�c;eX��,�B����=Ē��0	��P���9��Sd��_Zڨ(\�W~HR������K=�CRW'9g�(;ز�5���^*�[X�*h��Ə���lm$܍��ƅ����w��8��q*?I�bf#��
R6����ŕVT�XW>Oq5^I~=FA�v���CGnj�,��[���-���8
W�a^�F}/��z�MT�d��㕸�Z����OD�3����K�LF,N�9�
(t�o�'���Maˇ��-n�D�	�k�.�G�Ug_m`/>��v�)I:�$E�Qfއ;͆3�10ɝv���NZ&ݬb�QQ�i��i�d�S�{�	��&
'���ړX���@�J��U6��u:!�VYy1�����
���֥�q��|���o7�.�R���㶍�����p�T�St��Cn.����ȇ6���Ʉ����\��WJ� ��^�*)��e�����jGЕ�@��G�3N��{"��ݸ��ݟko>��|%�jw\��a26���l�7�s�J�6�]U(6Yi�:zݐ��/[ƺ�V��m��$�_P�NR�+���1$����~��8K}@��(���L�=�:Ÿ�FE��o��:��u��WD�B\�I�/1p�P��ipSnu��u#����Z�d�Fvj���ŵY�:�N�y�uG��|�j��=B>����$�mk��D��V�� ��[���4�;��'�h����#�� x����.̼��K�]U@#����vR*��.""R�RT�H]69%�5���$y`ʯ�����G%���^�/�7��rȰ��q҇�;99�:�^�e
�<{�ӱ5=��|T�%�p�`F*�ϩ��5�_�ܴu���!K�x��N�����L�Az�f	�n������_��o<d�&��[�y-�455˥qцN��>=��J&?�=���*>���+/+����-�3c��&�֪����s��E�v��l?3�k�PH׸o������(��c������z�C�$1ϩ�|�����2һ׼��{�4X�cu�A�ʜ�[v�:黎�mVn(��u40������H�uu�)㹄�� ��}.s�j�L���J-v{���ч����:y��os��-R��>ny�v͟>�*�U�ua�6G'7lYg���N��hP�]H�uU�v3�_	?���~L�k-zeU�A��ӽD�;3��"���	�*�	P\���x�pQ��f=��I=�mY����$qo��Ռ�̀��Y�n<���z�sdt"��dUԦbo��N�v�	^���&^o*6�ލ1�^�-����m_�����q�%-vzj?���j��ێ��IM13�_�u���s�-|uyhS������������F{8���Ƥ<�������=�?cވ>��yû�;m`m�u�qi�/���#Aq��kV����j��g\��7�ϱ��'2,GQ[gm����u�֓��2��x3�x2�ʆ���-�7n��AJ�%n�Qr&�ۑ������}/��Ctr<���K���/=E�V���?o�<�u���V���O�I����w�����E��ͼ���̕��=�� rvlل���蜦{6
�*_���]��ݳ�ؠ����I̸�����m$\8�~���&��e�Q�r�N�DҞp�-.u(�M�n��I�	��ڢ��`�ݜ�y�l$m��-�3�!�7ؿM�B�|vݎ��faeL����w/6���pr2.e7�۵������h쉼&sV5YH�b���X���K��#A������+b���;�(��!����n��Ι��:�7��&(�վ����%��îD����t��b�0)�t!�&mllB�k�g-����	�h;ym"=Τc}���{���bC��کjj�F:Ž�A�/��]b��Z�_պ족��D!'�s�U�L6�D��Pu���C��T
��d�K�/���:��������DH� ���5i't�f�4�
j�_�8_�L�9��Dr����L�b�~�'�z�)
���X�ʪ|���^�K����ָ52*��)	���0RڄN�ٻ
b�϶-��y����:���+N09m׌29�Pc����D���H�Wzhg�Wz�_�3�d%w���Ҫ!5��W���o����T�.�g�jRn[�PE�.t����iY���K^j�Ƅ7����s��� |岃��MTM��N�r\RU,�Bq
��IZ\����1ڪZ9.7J�R�J=�O>����這�C�4 �1���	�	�������:�Ie� �#�%�s�b�??�D(��h݌u�5(p��}���OYaQ��)
\5�'�0=�kd�1a:ame%.7��1�V(��Ԅ��P��j/���0eL��s$�Q�'x�@�|&-N������E�?ST� K�BKo��_��Q��ڐ����P����٭&A����{|(����5�m|�j6�'`X#�����>%V�CR��'�;��fAg@�p��t��ri�
�ͮ�^~���������IҒ���ȕzK�L@g�u��&;}���).|�ϑ�	%eeΨ�O��:;n���?%�2���,��&�m�)�7��R���D��"�}�4�QH/�"�p��+�x��6���}.��
&ٳ�������7L��Պq��i���˜@��$�g_�����L�M[GOq�	m�{����,4s���*Kb�o��/�(%�/-o����C/6�����ͪl��*�@7��dt���(���V��S�a�G^�Hlm.�Snm_������O 8f���[�����:ۿ��S��|��궷�b?D5��:�[�+�(���-��P�C���U��i��恱��E�~���Kl�)h���Ռ	��q��s�%?��R�2F�("�X�$����+�m�	 �+���L<:��uks}�xK���8�3���e/��ۅ|@WkS�i��Xp2$5[O+�����g�U{e�2��?���&3��)�I�h�du��]E^��'yau#��ln��he\S�#��<Ċf���7����'gʇuꆩ�;�57X�c��zM�,����:���V�S/ֆ��u�+Æ:���`�s̑=w�f¹�b 
���{�k�AH���	�4Y	
	�f_����<�vUa��'�����`
ϟ�O"�����Q0�v�6�� �8 �����u��*�!��ԝGQ�D�������.��Vsf���x�+,c����L�m�`��]Xm�]~���<��ْlP�S���T����EM(�j%r��9]Brr����/�#~9�{D8��U��0�*��l ���������I�JA�A.�YNql-�ې�������??\��i%pRr�W����"��PS�10�,9U�2�3�Z8���F���#,\�||ƼǾD.��N�ۃ��
>�ɹJ�J�pZ<\���(:�x�ȍ4�6�W���u4#^N�+2��.0�����\�-��+�l<E���$���c�ȇO|M��;�[RTD��\�ͽ��)�$
���t���O�K�c�Vs(���!���7π��7x���{��onڔ��46<��T]w¹��eEd�x���9Ӆ ��� ��yⓟ�����X����K^�ڼ�_���`q~x�r H���0�[���2�n*�|Մ�e�8c� Gm�Q��|ǃ&��Vd��w싱r��3>Q���}����͉<��9J��d?J�̛�A�,�ϔ/�����1�Ӛ.$#3s�'Y!�)�ZFb��2g���u�pa��ӛ������EW9��.�����.��v�e��K`�y2��}}}5�����T��7�W�HQ��j��@�3‧����i��� ����
~�����:��8���x�����9.VS<�~&|j����f��.�ȭ�L#޳�����$�ʮ�K�H� R��p ��we����Z����Rkgj6��O��~;��s$��,J�h����8J&���5滨��Y�§����]��Y�1�1�3����p鯿�Zq���KIu��^q��S��&�%�nLHH��>�?�ArQ�!R57�Q2���M��Pu��w='��x겇 ��a�������`��6� ��7d�ڄ���!��aZ�)u��jA�=��$$�'&�����@�&2mK��h�0��P��Hm��[�H9쵃��N�;e�ϡ����7k��`��!�r�w�D`�S�S��Ԟ�������a�d]����eLXYp��D��P����4L_�
 <÷:MJ��\v�nqE��1�Ǎ�ޒ�hfWb�	K䧝���t9�ʏnen�)��L�R' ��;����;�]Cè9���H��SKk9B�k��ݺ��|c쉰O�b,�ߝ��8�z�2����+�I�U{��M��\���)/S�ou6mU��:���¼�a��n-pR?�Sy�
GJ�Ebd��ZA��&R,�������Q��ĵ�/�
R�s����+ks)��/���:�?�Ҭ:^x3�S�<o�A�C��2��������{V�{�M-��4[����u_L9�qq7Ƒ3|�'m�`�2�}]賓%~�Xru	��>�9%�y* )A���������ǐ�1���]#)tk���>CU}���~�Q�x����b�5����2����3��o��5���J���g���ůt1Rt�,�l�1gᙳp��:u��?�)�[w e7�W����hjjB:(/�Q\���� 57�KjP�?�yb$��ai\q�r���̝(�<���� ������#Z�e���Mf�Oc�@���<��� ��ϕف�ԏ�l�R�(;?��k�۶�Q��!�b,'N��^�|m�?��S6���T�������b���0U'#�� �#�no����_�G��iUM�Zm��ˋ�9���VC��4u���i����lQב�����L^�Sg�k�V����լ,��m����E<p�E��e_ӺT:?=P��~m_B�L��W9�<is�+U�Z�<v�L��dʰӞ�q�c"���Zw��5P�w=�z����:�����w7	hF���~<D`�dChh�yc�S�4�N�(�u����,&��{�v��Ё��'�n�esi�8���� ��Q�|ß3q��$���a��B4�	 HG��O���ku��:^j��K�,��i���m�����AZ�����W�1�4�/e���6��S�|��}A*�6��ތMq�B�K�ē����z:>�l�d�"�zV幚T
�e1R��������l��S.���\ް(Q��k��X^^~=J����`�M���e�L�9���7�4�<�#G^[�Tm���y�w�K�0Ĭ!�Mԏ�C��t�:��~&����F���kN�W��,�{j�X�Bvz�=nO�^l�2O/���.��t9
�۲D>�9>�]�����hsH���%v��V�݌��-c�?h�}��h�
�B[��<�������c�AcA÷-jek��"�p=�A������64����V��|2s�A�s.�旑E��js붖nK��f��?�=Vȉ�C���)ᴸb:��J(�W�9��|Hh���4�!%�p��ʰ�B#-B*5����=�_�{qq��.{�H�����X�������/���5��%�������K�5֗��~H�խ�yl�-�3��>�a�H抃�C_O�~��ˠ��arP2A
3�V���@���&���:�K�x�����E_�_L�a�zU`�_F��+���8����k��5^�:���($�N]&����SI��� U�j�±�k��h��J!�66�Ї��M�	�8�} �O��ϟ���kg�i  0�_��n���l�˰�����k)۫̄�m��?���.�ޅ>s�a�E�M�co���**^3}B;�\�G
|~uZZZ���˛ߨ��͞�=�[��h�K*�N�qb~�����@Tᦣ���
�W�e#i�ND=��\c��GK��7�<ǚcΙzx3��'�hqY�A������Z\铓v'C\��3���9՝��%E�3��i��Z3[�#��-�;��D�&�|___,a1b�DB��\��u�~��T��d23E����9	Kn��c��%�N�n/��VU��k�Y�k��(Ґ`�%U,��)�鵅c���=��R�P �G4�;�۽�+�Y��[��~u���Ի�\;]��]��v��U%14����Ǩ�y��	b�뭭�ϖ2V�vd(�>2���.¸ۿ�J��UZ�ײ�@����C��)~��{.��g׽���sT�����UU0o�?��8�_�Z����UnQ�LNN�MǧO;&K&��/h�YWV6������E��Y��G�e�B$���zn���K���l�<o�CF�P;1�U����yK"���<�,�<Fd-E4�i� ��Y�j�� \ԏ>���ٱ��x��u{{��~��B&�{hԙJ��ȕ�ohU}� D��?t9o�Q6�rii>��r���/�qg��v�Ѝ5�������U$�b�Kf�|�(�x%���w�>66
�?��/�"�v�yϯ��de��2�е%��@���qr���$F5�1	z1[����e�]]���ʪ�����֜ԏ8�(��~� ���sysK����&SJ[�SYvv���]�x���s(�U�����?����n�Q��by�>5'�+��?aaa��9P���Z[[�R�8���V�6��CR$�_��tEKQ�S���`��e��A���s� 3���c��|@�/�QD7{�ױ�7�eL�ϯ�����E�{���`����ٙ�4��,�m�k+�}ܧƤ������dFƟ�����uy�min�SYd���4�͝��;�\�#�@9��W{�:`�zx�Wo1��վ{��Nx�M`K��0��z�uȚb��~;U�:��G����y�>�y�A�8P���ۋ�l��6Ŝ��G�� EEEe(̡��Qu��畼?ޕFu5�.Cm$f@KEb]��I��nC��/I�]���ᜉ�	��^��111`��ri �H7~�d���KY�:%������7IY��ĵ�$���9�Ž]Q
�Lz@��y��R���
��w�WDcZ�K�~kk��sR���T��(��2��WVZ�U�p�ޗ�0O�R����YJ�h@���oj���WR���YY�����)0���ͥw���S��a�sW��(�=Ĝĺ�+��:;9b���MV���瀨�)��������u�I8�I�s�֠4�ځ]����xJ��skj����0���Z�^@�o��;�"pl02x�-�gve-88gZ�f�~����/2�ɉ�\NLLLPH�Z���.6��i�M zK<-�:����s������Z����=�7R<F��A,���IO��a"CjL"��E�R)p�����#p�YB�j�}��{�h���!�G /X؈KU��vB���Av�9W�g��uujri4�����^GaH}x�&�����Ǐ�}�� ��G�C�A�xΪ���ru[U�l��'[3.�>]7\�Ǔ����u�>��������`��T������|�9	�{z��M'�N��\N�|E����%�1�'�)��f��/�Qx�tϔ`R���MĊ��w�~Lm�f�+5��CĊ�l��*�mi�S�e�I*X���r�8k}Y����p�p5��sݦ�O���M�%���|��+�}}�<���X��g�uPH�6�'�أ����g�w���y���o�Wh� �����|^�6�¡�������k�4'�$"�b�X���<������9�g�����]Z�=0�lR�^+A(%�,�]��_j�_�{�Ճ�j��~>>�h������*����AyF�ܺ�Z��u&���SQq�|�r���3$5���Y���3��n��� �������6b# ��1�G|w���� U��= دP�;��s�.�L��.��M���ʻo�(�Cg�� �T��L�yS��@�|�'�~7��`��Aon`��wȐ	@wM���ߒ0(s<Iذc$���.*ػ��Ƥ ������%�2�F��`�-	�A�~��j��3�������%u��[	H'��s�a�ڵ�f�9�,G��i����i����>�ַwpЄ2����X�a

B�댸Ujik�Ր�7p!� ���m�:?]�]
<\[k�ض[�����O���v�f�jVu�a��G��� �p[@Ʀ��aH�'�#�}H	*l��?�*�+RZ��9���-������ʱ��?o����YS�u @��z��j������A�h	:��*�[3�o7�(c\L�59��>|XV�A;���2p��2a���U�M���A�o&o<�.�pd?\��n��ek52��1B0��)��p������q�B�;�Vj�ف,��fe(P'Ooog��#��?W��ϟW�8�v�ߴ4⍃���(�|E��[���ְ N2���(>�?&a�f��Dt����Ç��zMJ��	#��oIpqsG��W���&cX�~��գĞ%�E�{
�A"zx|&��������cccP�_���]@k�1som���Vr��x㦋���kk�Nõƀ��H�f���#�`᪕!?P���%p�����8+�:�ekvv�h�Le��^�g�k��P.2�ձM���90�wΰ�"�Y"t\�Fy�w�����@�w��̴�p���h�^	�(�� :���f�&&�&������naq�X��N��/n:
.:
�5Ӟ-EZ��و���4_"�8Z��#�)����+��g��@�C�l]Z*<( �2F��e�/�{�N���q�*����7p��<m�t�D!�o54���k�wq!��YU=謭��Z $±c� �3�n���~p �M�:?�z�bY*�Mcf����rn�h	{���%j���89wv��5xh��W����y���������q��Ou�5g��!ii(��S���3��/�9�5�J#�/⣍��!�31u���>r�C��ݣ?yR�=�<��P�R���\�w) ��^(p�����2���9~���t�.Dc	^�щ!�=zgz0�8\3�v�Y��u*�����9A�}39�8�ר�Em�j�nnnNMOR��Y���mh�[U%���M[����kG��n�9hkU��`q^YI�#�%>�S�ҫ��Zr���
����g�D	�|���g�޷o�ǟ_��KKY����_�4�sRG��ۻ�����ghz9'?_�['����ܝ==Y�-��[8d���Y�?�X��Ç=㗑?����S�;~0���7��,�>����أ�:�L�2B=I*����ZO��������U��oy�2�Uɮ.�)�$��Ii��CKa��� �Ǿ����
rgsw)�"{:Y^]�s*ZL\\�9Ǐ+�І��6� ��0���G�}a�c+��˶���SSS�SCP��"`
v���ay<��!K$����fp��&JVb:ğ�B�B���Ag>)L�w���� �������'/�xH�4��Y(��便Bl�TK`�h��:��*��X�i�|FF3p�������q�|����*-��b�J��|} 'Q��號bd<�o��ȷ����]����;Q������i�!&h/:��Ǭ�J��ݞ&���:�Os��f�?!!��DDr�I0X7�$B<c���n鹼��%E��Q�AL�2��*�S��zϗ#�����:B�7��>Wɤ?u�s�U�e�7�����F��o�^^^^��yS�=}��ȋ��xZ������� ق��*I��yH`.=B���'�,�r���D{����ث��Ej|KK6}����Ȏ"몠X����0U�$ǌ��޶7��+�"&ְ<'#����K�������Ի�C����)�*t�D �h���9PM�ܪ3�va(���f*݃��7E���t�Vx6<��������;���j'�;�p8�m����ϐ�JSGL�򅱒t��U��NN1���4Kl�q����$I?HUnG$�Jؚ�x@�e��^�`��u��=`,�7�\��6?[��!�E������{���t��4`X ���!�<�NS�~uV��+��W��d��Q�̭�P��/����� kD�%?��ohٶ%k��F�$��kf������ཽ�s�TWn�E�A!!��o7��yf	��Ş�k���v��҄��3~>�Ga�,�DaD�U2q�j�b>���Ô�\��<�Natx�J�k�"�]]]�..��o�����":���~t��ڒHJ\!?91��*9tgUV�ࡀ�FE9��(����(���5��������H4`G�`�����C�[�h���X���a:EV��ϭ�-0��{����'��v�:�H��hiI�pcHJ��Ȗ�N.��Y�����Mԏ�O�q�n)*�_u���9��� ��0:�IM̌�#��F�����L�jռ�G�s��aSH����4�ݍi���@���o�.L=�����^ r4�����έ8,Ouӎj h�g��߿�]�a���rre)G{;;u&y�g�7�=��|
�n�ۛ�h��''�����V+I����?[�����$����Yp���Х&}q��;F�y* I0ߏ���d���Ǵw�.��c=�A����E��[�q=]CM�1K�A�߰����ʃ���Н׾�<]�:*�����a���J �	��'����y������9<(��FJ�6wK�����F?��]�S�-� �7X� 3F!�i��L�ݹt	#��w�''=PU����B��EK++�puH6PC�xL�km{\z�c��]/�#�]DY<3\g��gF���#���u����3?>�sEuZ����s��[[�E���Ԋ��0z�m�P��P��}��J������eX�������bԷY����,c���"Q}a	z�҈�1kB� r��M������A��� �6D Z��\�H�Uշ�04��?�ԦV�81�ʖ1of*�7S�M
t�fw.��_��)�el�mM������,�($j�	��Qƞ��ݭ��a��K��1A����kʘ�Z#�v�cd�WQ��O�"D���,
ʰ�BK(��&^m�f(�����v�c�/0v�����ۺ���g�ߑ̺�����|�7�09��]!��LPkOd�#j��D��	��A�*�/�9L�ǙX���A��/�3��)':�"g53�KKˏ-��F*�d����Ff��ؚkT�&��ֻh�D>��7����>��8���ȣ5[k�hyճ���6E� ��>�6(��ԑ犿�e��=5�3�9�����f���X�]IA���C0����_�@�A\����e-z	����/Q��� �|$����:��+W�i\ �uMok��k&E�=�7Q��ϋ5���`��i����~.��&��f�w����>�\E�Oz�z;�.�e&��V�j����oq��G5ѰWkz�cx��|v.�>��H��[�2O�ݽXk`-�*�� �֝�Nr1��!�'��?7(s�Gqk\��Is��CL{�1�x�a�Z���ZP�a�w�/���h�q��m��}qt���e�������j�`�p���+J�fDVm����p�n�	(�0�����ç��.b,ht.����7UPb��[�{Ṣ��䄺@�N}�-EJ������`�h�6�K�v�DV~~7��[�	@�ܤ !�+x���]�w���u�&K��@����ۅ��ۻ��8�r�@_��b�ȇ�	�i��nG(_mV�p@�߃��8���C��]Bc֔��%p��E�H��t%�_�e�AO��o�{N��P1�E/6iq�ߒȇ"�*��g��7&slQ}��R�#�� �E<�GHJ*�-�G�W�R��^G(?�C5~]CC_��1������+o.��u��6��ǀ�K{�����41�����:K$�X��M�� ����t������5&��d D�)��CA�P�����Ѧ1��8W����i�hU���ap�-�������|��]�or삂���W���v@��ywJ2�|�W�, �6����l������C�@h����c�n�����}���@��j�,����N'�)���{����Ԗ�Vj��
��<t$�Y��_��x������B���H@h���MQ����~���!�;��O�m���%��<_X�9�"�!F�zD?6��u4��S`�$F��F���(�fc����4�d�����h+�P�'EQ >���#�� ��A�P?�I��eU c�{.�.����#������B�^kq鴙��V�JKK[[.�B����S�l_3w{�1�ԉ�J!�P�t{�v_���0`ǨW=x{ep�1z�y�T������n?�����&h[�pXt] �h�I�$S�pKKK)<(['�{kO���/�)굹�-���";���d���2�~��~(#�3 �zP'�	h7�\\ 9�����ugT� >��Y̨�3��`҆lz��*2{
F�dU�ߛ��	�.���l�u��r��b��
@#��
����D�)����\k�H
��MF����u}hEjf�&�v�[�A�� ����E���0�=/'G�y��|��P�秈F���+M��s����ǏOe>��g�F{�� �e�F��(1��B-�|�\��!������!MU9��{{����������l�\7�|�+gaD�2ꐉT
�¥li'�<�2�6*�e	�-1��F�7N�ҁ ��qvg.B��J�aI�a%ǼX�1x;�m�7MF	�X$&ϝ;0-��6}p���!��X�q�-c�]/�؛���53��w�Y�T�h��s�\����U]@�:+���j�T�<�QM���9�����
��)m�j� ?�z�w	qR/�&��^���,��_�T��S�4�
�F!( ��6�9� �ޠ�@?��|2���P}��J$, �;/,�uV5��\�0�?qҭr�7�l�Rs�Jhf���n.U,���)����Iw������*M��������+uۛUc��
�����#�����_��Ä��Q����~���7*��p��%��7M��b���^�rJ..����H�������(�"�����ꘑ,-� p�U�f+�i2(WUs�����1f_��yxyM��&��Nr`:A$-��4j��a�Kp#�Z� n|e%p� x��8�{�s9jm*�s�!���7���y�H�q��HzUj��`�az�+�C���ZÄT6f�Ez�,��|�ׯfb1��.
C##/���@<�x�`Y�#µ$�$�_adc����ը�ӧ����j��lS�t�V��#�}46��ꦁ���3����(��E4���glчQ��%��IU!4mE�cS�[b�B;������%)�$wb���m.dT練IU�F��4�C�;Qxٞ��lm�(d���+��W,٣8�3�V-c�d@NqVT�^I��=��+F�x�|XlH�|�T�m���Kx���1��?�.xr��]@�*�$ IV{�r�3:�k�ϸ�~7�\5`!�_ -�z`����������S�&���O�F���+���c?wa\�m3!R�/����
jH6�ps�oxbD̀|��UUU��fz(F"#n��r/�N��!Cfac��>+����L�aG���/��U�a���Ч17r���(� �s�ږ?6h%���1)�?�1�U�WG)	+��+�����G�2��2q�[����m��
�1�q췿KQ�Ԍ#�s��~�� :� I�=�7���Y��2�7�.�9����d��p�7R��М�F��y��@�o\"�r7&�쓤��e9
���}������P�Wi��%����4�f�b;Hߵ	y�3� �Fh��GtF,����W�(v0��޹|:�z�}������188853��C�	!3��I��9@�y��;��IG�ST���[�����`%y�/Z,hZ��NM� ��~ q�s�u=�+�l��5 ?�9iiW���#hB���?tvuM���VQ��,<,<|jidBW�^�+�k���x%�*���Eg�3yB��9�]V��:+���䐆P�(L�ʻ�����ZTPD�i�fl����O��h\�pL ����{��ҁ�{�o�����e�Y;�3��L!�G���&_2�燆T�ˬ�`oN^jΡ�T��x��"�E��Ў�D@;��^���^�RK�TMD��àD��1o\		�b��ξ���h;���r^�Z	�D�A���I�L|}�
!nA���\��!ڛ�����[4��W� �K����A�L�n����m��<,]]]�#w�;;:,�1�@k�x��F��~�nD�Х�߷$�T�B��<ף��0@��k�g�*��+���M83��XF� �e#޸�w����JlZ靆�Zs�h<۹�Ś�R��HIؚ�(�5aɼ���%cE���!�U�%Y��h�{�p)[��B@ݰ�7�����jHH�S�B�c�%�4Hj��LN��Tf�7Œ���(=>�]b�c���zF�ӈ�E�3�Ä{*ʈ2t�-������H�4�z���Z�.W���ʰ�-Jo����&3�U�}�����%(�ă-�"��i�*́�\0�T����=EO_����8mF+&&��Ƽy-�|��.דQ�>tB�s"p����@4� �� ��c}�|zk}.��7~�r��VRQ��X]�����<h��Rmcn	���KK�K�*�1-c?7{0�*D�x�ҥ����]K�H��@7�@H$�/\G�	�ߛ������堼�?[@
?;$�Kz'�I�bCĪ���_�ҹ		����?@�9��q�D�B��Zً^bI��C��Z�����D�:NNX����y���0/fg���Q�����<��$2K6�y�Ə���N�����<~�?ʼ]���:A��mCx�|C(�S�/˙2�V	E��:�ќ�Z�L'@P:�u���)(�k���x� ��cn��!��&�UU����׫�S�R�/�{����'�k�Y� I�֙)ņ(0a8A�JH���a**#�ZY����$J���IEa�"Zx��XE[;���k� � �*���}3GV]����<�1��04[1J)�Oef��,*���EzffD�~jCb
�kN��/����u��� 4A&=|M"�!reW��59�a�:��hE[�3q�f�Yp��Q����������^SU�i���
m��b�DY	�2��8裷1h�֮�������H}���gO0�*�ٳ�PSR�;:���̱}��}��� ��`�;�\ �����wq��/ ,��^WW6PA-�,��O׉�R	;%�iv�
�4ik2a�<��k_x�I���EX�z���:z���+�ߒ��Ё��F�C�m�3jM7>uz�|������������|*�!�=0Ѩ�b�NOF�Fx�)�ٖs��[?T�U� x��Mc�/g\�'!�WOq鶕Z<�ScBL��
��vu4i��u��1�:Z��#�n]�e.��QҠs\��Sªe�0����G9`�3^đ�:���e;����%�To��c%�2�QR(�Ch�"�<��)�H�2��IHu��d�L�#!eH�B2d.Q���C��߿ǽO�:gkx׻�^{o��n~>��d ʮ��u�� �&�����`0����u6__�=B1�>��2\k����v�����p�@D:Gj�oŮ�گ��|(2�2��7߾=����'�"�e�A�I�K��@�Y�����`�qf�YY�Cʱ��i\~��&�_1o��Q�t������\��_����{䨪�<�QDx���ȿNnT ±L����6��?ξ��k�(:��^�j�Z�Z��H�~�9	�����9�~O $���}���š|7X��Fz����>'�yc�b>�)[�����]w����pt~�/��?�E��|��n]�n~QӏO&
�(w�C0<,Xq������\�"tk^9Gc��e]��{��B�/1�va���x�oh;�7L���ϯ�a�{qm=�3�Pm��`g�|� �2�8:�y��O��1��E�8�2���_s.����1�\ �~{�{������WRi-��;�O�� �*=,C/Ni;��j�y'��߽Gߜ�T�4X�� ����\��~����?ο�~~T�oq�o Xஞ?Z������l�-�]��Mk���6\�Yl���-�/`��¡��v"��z/�+���1^�u�!�r��	��3��(Zs��,�0�rL�=��-�j{��u6��y6Pd���f����$�g�C��J��>�+~�C~zE�i�w?�~��º�#G9o
(m	:�2=��ȥ��3����Ą��rS8��Eb�R�6��M/�_�_��і�Q���x�Q@�qq*+W��vÎ�1n�;#w�Uε���������r�^j��a�!�5��=З�dR�ҥQ��ĝ`��A
(���� ��I֊�.n�ԋt+r����[�XPH��+w� @��#~oU9�	���4���r=<,,�I�p����M��׿[_w��n�=�z��b��#u��#�m�_��f+/�	{.���ayG`mO�����&�e���U�M]����GTT0(m2���jd�H�,m=�R8��0�� ��|�9/�r�i��v��{��&#���a�^����c��=Ƶ�cƖ�%Me�l ��!�3e��5��SЊ���T�Q�\ �����Q��!��bCu��̻��¹�/l�����:���he2�2�x�7+�GQ,�����\��|ZȔ���_`���7���9�+�:r����ߖ�"�]����Q�yY����q##�OȽI+u�v~�6����G [�^x���X��p��-��m��{���z{<8�p��sO� ����������p����B1d, ��0�*@��ó_��f�@��4?�V�qz%IU͍���j�`oi94 &���D����RG��|1�X��.*�@/a1�m�D���eהk�$覴)����b^)[/�:���n��(�������#���
�Pz�Gutt4��6t��?���yS��&��2F���� ���ϟ?ҹI2��U���C*1�&?�/?��B_-n}t�-y9�,N+m���:Y��Zt�`��&x_Z�������P�U><\)���*������9B6<i���^XT��It�M�����`��G�_��{������s�]ʡ`��X�ƃ�ې��~6�6U���������v�����|b�tXm���h�6Mk뎴7i�e�1�_'s���������
�>^v!ݼ�av�!D�
H&�:?S��Ӄ4�OB�K��z�'H��]{����fF��+�Ph�z_�C�d]n2A�__��W�j{�h��8�"��r�o�����}A��3��Q��m�6l��7 �p�/��'�]�g�a�em���n���Y��{l��yI�0o�}��̸��&���o�kd�U�`����E�wYVF��b�g���싘��j�*߾�1�KdR�D0���e�_����:t��r*_��Ҽt���ކ,��o743���Դ�W����P��@���W��� L<��G�.�&'���	"�p(�?J0���@t�	d,�?��+Cr"|�a$�BƤ�8��ɚ�ˆ���p�ݗw��Y4jjk?{�����i�v��ޟ�x7y<�,�E�m�Y�O�6,�/y#˕=�Z���n�|�BB����.����ĉ�0Pp�-`6�:KB��7:�~<��ڟjQ������"}!�ئ�7T�5Y"���
	�M9�M扺 ^լaa�T��o8��M/،T��w���놆2�y'䖵��c&�,N&^��-W��M��*�q�+m|l`�u�ǏG�u��J066�����%d<��2;����nA�ϐ��ٔ�LF��#�ƪ�� ;��@,ܻ3�
��5x��K�`*�m�����4���32R�&|� W�t���܄D�6�g		���Y��#�4#�:]����lxvGv�����*��Pů�eN]j��/�~B�u(�����9�D�l6�khkG��jI[��x�L��f`]7�I.�����p~o�������6-��X>k�Һz/�8�YE�ӧ��c��4�͔2�<��]���ǚ�����~L4J��
�r�Hw�H���X[��q���T<�ܐ�Pfr|���(���{#cno�s��;&�n�wr�������*�z����N�AѵL;_�8�������Fr&o��Vsf�ǥ��_��ʲ��Ns���*�Bׅ�~]�/�tL�������d։���B�v�7AWrr�w�z�GeUՓ���@�jsv��p������l�H.�9j�j��t�=`����A�w �p�T�u��H6����p|����^z?���O�t�k_�Z*�:9��ɉ��5ww��9�ZL1�J;�
2�����艺o��z(��'_^� �p�4x�*������s~w��F�P��!�d:��G�M�����¯�]w�J��B01�����"1��&$�z�����6(�Ι~�S˛x4�(�������79�̴o��Pr�
��g�{�%�M��rĐ k/E�{�#\ggh�j�g�iQ7.��5��kn缩'@�|llL��`����"�@G�ɜW�Ź2���E&�MK�M��?��:�����A}�'~�;�I`��R������h;��{R���888t�?����^���ɱ�ɾ`�9jjiu���E,�������x|����rSM��Ǜ��k���e'K�P�L��y.�0^�U,P���j�U�����ɜ�Ef�N�v8+���n�[L��)+���p}�js�l�R�����C7zHQUՏS��)�����+B2�i��T$�� �=��UP���*��+
j-�Jz�v)�wl�������b��>�X��׮��ݵt�>�w}�a�9�5�)�1�eÆ}��K+ǆn�q���2��[2�&�#VC|۳�=t�Л���A����2j�j���6ۏ���]#�c�0)V�2|���Fp֔����,?'��ԏ����1ժ�~E5��Ɇ	��?�	4�2����}�`��T�|}}G��'�����(�'{!y���F��Z�j�,X O�O _��Eb���	Vk�D��8َ����1R���bd��e��w�T�ģ`XR������g�T�P�}$fQ��nk�@���j������h�		5�j��#���/�p���M<����Yk�yv��%R�n%�g���U���ޑ�����)��(���2|��]�T���T��ѭ��Ј��\B6䓊t�#1����[9!�c�&Mf���ڴ�IN��-<���t��󜤶J�l�xSW��u��k:t���V��F�K�n#1��߾}���s��#p��t��X�_��ű�~��:K��&.�S[�G�jq	���� p��T�v<������G]��k�l1�63��U�d��6^J�)&��b�הzQ?x�#���ֵ	Z {������3�f���D	II�H.J�K�5�?��*a^L=��!oN#7k	���M �p��,xeޒ�/N_�$�G3���iڴ����WQcc.n����������}�f���@��ޗ�'���{�]@��A��=���˛uɚ8�N�������K��`��|�B?�X,a�׸qe�-}��*��j�����)�	snY ����=�s���W�+�5c�P>4��[ׯ�r�W[]�{�#ŚF�����V,�8�[D*X��9H���ɡ�U�l�:�>���������������g��}ddd������
P���-x'�=	�`�CG���cV#������ݧA�:^ �e��`��K��5d�		)ӯ3<p�S�����g��;LZ��� Y]m6g�w�y��%���nZ�p�YCPx��� �����"��=�@&TƦ��G�eFD�{�y���Zy#���1��n4���=��Ku��F~�OƝ�9W�w��~qJ3-Z�î����/پ|�Y��	�Dq�����[�frVX��5��C�y��O���]����n_��v��]]]5<
&J��B^:���u��Z��$�L���|���{2N	�rh��ƲiP�R|a�"�����@ ��V�]��ȹ��R7:�?�a���ۛd}g|tT	�5��ԏՃ��ѵ�U����V$�g��`���4�
* V�y��3o������q�_B��whA�'<n��Ө��v��K&��#�*H,\M^��F���;{�g�$k��>\
�s㤢5�ߊ�5�{m����>��>�N�Ie9'��&��U)��E���#����3T��o��]Z��o�G��nDMH$.�9�?��i��2��\�p�H� ��y�y�*ס��5<�0�������1.��ц�@D�]�+�����6�����h��x>�F����O@Nl�Ui�4-X��3�^^�]�^GXL:�u���X)�4ɕ4��/|O)�O*H!���k�b��[#=��[H�}����emR~s���N�R���#���='w�.�'��4�w��D�����]"�����"y4>r(�k�����$��E\�		g�j���Y
������B����_��𥿽ie�WXX��yi=jB���Q�@����V	��9�� �l���0������'%���x��#��> ٳ�b�aӏ������u����8�<S-+��j������ey,�y|�k�f�!���\BB���`m���u��c�]- �C�ŧ(/]�x�cﬅ������-JR����a�=֗��j �;���Ѫ��n8�.u��ߥ�8TF�K]]B[��'���V��.���W��z+�}b�����B[���K��ן���KKK#.iij��^Y���P�5��OS�ֳ70��c	����ۮ`ۊ���Aaa��˱����{�V�M�5<s�A�z���_����t�O�������p)��;!<� V�P�<�'^?���%k��ȑ��uN��l	��V3����g�"�H��2Ӧ�6�U��C�?�v)�;�):R{6������X`\�4#���U&���&�8��s7Y��ϒ����Սq Nv�r	UF(�"6���h��>.[|�#��R7�b 0�K�ܼ���|1Xb��$99�y'/9��/xxP�~v���7��ߗ��_�!ر��� �^GȦ�/	�8'F@�7iD��h7����c����F�%V16��D?Ö:�ɇv��}��gz h!YYY�8�xr	��'Q��A0�81
���3�q��ڼ5ܷ^@��%��[�"�(^h �8W߹zI'=��d̩�$H�0����_p�ׯ_0l�7���m"��R��X�7xpX[Z"+��l��p���q����l��H��ƾ�Cy�쀛������27��wCI6��[��b$G;t�uyrŴ���&D��`��CDt��2���DF�_���`t� ��������IwVZ�QQ��u�^��AgXH�蛬�G�D�!w�n��������	��3����}��$���M��}����%��?K�0����w�Un��ԑ�.w�0�~<��̏�4��]	ET��cX���X`cҰ��(qXY9�v��#���g�%?#��� �a �n�÷����XƷ��� ��IE�MHa7����n<$-l�dݯ���/�:���DA���=����g;���Z�u��E&[���V'�8Sm�D˭�؁�`�NuC�������)���y;i��KǛmR(�6.�Z0Ȑ!���Ԕ�\Ν1�inum1b�Н� +w@S���~�`���С�����*f�o�_ ������ݳ�Ȃ9���<u�N�"�X�����'j�l�v� � D�3+��	��+H�(���kK�k'�Q<,�OS�&67FI3FJ��9�b	�|#~�Q���AT��e�B`�׀w��g���!�PH|������L]��뎬>˳v0w���.	���C��� |��0pi�b4\5߹���(hC;�RL�$'��9i���L���L�p�DP� 2�s'HK�gnB��Í㞆,���s�G����YDs�D�v<%Vq��+@;e��G�M鄼��""�\��g�X��=WX���i/^�H	ω�Cx��c�u=�:ܲ��q���h~O��m��XOJ_) r
[8�	ȰZ���_*lNe�jR`u����v���`���k���2Q.Cd01][[��U4S�p���X�h���i�w�$��t��UR�2�yP�#�l�F�r�yv g0��Y�mZ~b��j�����>��lf����F���j�C��2`N�[BU���G��.~�������5�D�E�ߗ�{�Ҭ�GJ���?���2�P��2	��{عO�29��J��K�.���r�+>y�R�&pA��Õ�h���o޼�O��
���ڪ�7m�'�����b5<��Q�}Q##��
��M��
�� E�X	�Nr���̑���&�y $S�����3�}<��˗�%GBw���ɂ!�K�����@���������'���7
�c[ed�pKi�ȏ}�;j���aR~���HC����i�Q4b~b�G�}+q�O��_]�S)�~�Y������֡7ϴb�jj�g���Ǔ��	�V������0� +�.H��s��0��l�J��<�;6Q����%n}L���~Uy��]�Њ�֛b�)>���.�7����V��j��$�22�$&��n��H��8@Ӵ�L]�hUjr��
6ρ/?�t������&�n�5!����m�c��_�׳��v=��߿���"�)���J�5iZlx%=}W�^J!)�
2M$}�M���E�+�����&dd� �0N��|��B��ӳ��,��/��iffV�C�Mț�:��:_�ĉG�E�%͢�C�g��ӗ%fER���p�3��G��Y��%���,�?Sx�"��`�f�փ?����ſM�CDV���`���0'Q�E�cz���㫿��T�hhh��i�.�K*���}M[������o;%����m��pVٸ���Q:70�¼Yl1����� ���g��c V�x��<o̴���i[��2B��C���Ϗz�V�$��OF��e�3�9w<	YS�=�2U����|�lJ=�y*�71�1~��72:��sr������ѩ�1t;��#s>���]�87���oV  w�!�+���(�f���Z�RF9xuﺶ�l^ o<p�ӑ�I`EK�qi��.7�,>E
��I�F!VB��{[��֋vE��d����5��x؁7:�.�x�0P7�Q��˗x�8�Ltٴ]���F�Oj�)E^�/�9׬Y�I���	�_���G���2���`R>~��~���y9��MC�3g���l6/�_�b��mp�	-#��}����OX�RQq�zb���?@��C�-P��4��:������iȬ ����M�r�[��b�-�F>4�%�@��&�v1�犾����Z>*������~�� X��=���)7�v���������n��o+�ș�^�Z_oM=qW���ǉ5�H�Uyt�-�IA�>�>B__�G}LK:5�̹M�! tOO_��ˌ=��eۻ����Eݥ
@��<��5�u��ub-�T	�B����x�=55<&
#�Rd1���
�i��JBN��0`[�͢^J.$]������(xCn��9�:̇�+D>i�ֵ�T)��y�Y{i:�y����ԅA/�V���I�K���d3�]}xs���C)�ׯ�|�soI�o }���� sC�+;�N�B�OO�� #������[@�h4��:����dރ�: }w�|�se �e��zhL���!���X�t�ҥm�� ��Ӭ���jj�D�����\^��Y~���L���Ԁ�H�8��ׄ�6 o�$i��Ջ��q�s����$9N6O���Ҷ�������������<����wG��ځ�� X޽6Z���Gÿ�|!�f�q���]Gbb�y��GU�4���Ŧȏ��wT|���~��� d��D�5A\�g��V�gu�����6��>%%%�E;33�Eܐ��?c��H{j�,�"c��ͧ��{鿅?�,>^KO/��4 ���S�!��].$��}&�KAwvԙF)ρ�K���Z<i��;�k��"4�����Aj9��X���k��sg��[�f�e=�O�EI�x��9#�x��F��۹��S���OLO�nkk��g�/���<�o`�D����Yk`�*⫴pה��~�Xё���ӬC�/�,;u/�� �gΗ������ƅ���%�&��a܄��@��w΁ �޽;\]S3&��x��A������MP+�o���:}�	 ��74�Lc��Ç�{a�sO�����i�����=��-W��t�}�(��!�ce%�37���\�WcX)�/��;26%-�4 >>P �T�rz�������x�!l�����Ss�˚��M_� �Ά0���Ξ?}� ��,6��i���U���NH���(�Wd�n��� �&iZh[��*�V�Ķ��ŋL��hoN�)	&#�2�k'Տ�7-���3K=>&���Ke��v��%�	�K:�[�bKEm�R���M���n�o�=����?>9�J��$�my�������iI�A������}e��
S��R�E�w�� �u����G}F9i�����"F6T��rhh(���wIH�� ����R��b�r�.�>S|��`�%�R(����݃37 �m[P	�ھ}W�'�z����P|{���F�OD�G ِ��HL�E�����p��8�$����Iv�)�3��H�,OǤ2����pIl����"a����C��N`\Dث�}}*`�M����;��׀�������������Íۍ����(I�!.G��hL	�`�QDI�m{G�Z$ԗ����9�ӴӦ>�����a�_k��R�@h`鎌��T�@�"0�������+^�)�潸Q�ބ!<OK_��d�]�O�N/y�h��O�t�O���ˊ}�K���q�΂��,"���=5#��k��U-���N���*GV~/���?s'sM�`ֱ��^���\�깐�׹�x50.�0Q~�3#�&���v�`:h7D@��Ǐ�.Z�$ X�0?�Y6���54.�i���V�^=gI�� �?}��|�x��*�w$&)y����=���###�E���v��<�v��6_E[����P�?AF�ٲ�a ���S��=HMo��E����]�B`A��f��u��=z��s�mii۟�F��T	<��1|���8;�XT�����HC���f�wgg�z�H��7,S�O?�^&�4�ge{�����/y�s��u��i�sg��^�L�#0�C#}�K �c�R~��e�"#�*����[��k�瀯!�R�A��Α�D`¨`C�7/�SE�|��W��(�����{&��<r���R9'}�����2-6�u�2�>\l�K���b#sY�� f�VF#^=o'�'H'�*�9��n�Ց���a�Ϸ?c�O�q��*�#S�������^F}���#h׺����K�g�P&CO�0�:r>�ii1qq%�Zb�����kJ3;uʲЇ|y% pPv<j:��
�f��m�ٗW�#X�a������ů��1m�SX��9̲9�Ep��*�]�:��<�Q'W��=7�pd$���;�DcHKK�	 VU|��sC�,�4T��Ĕy���P�X���f�Lu!���)y!��S��l���O��� �F� �� 	�Ωz8�����Ga��(
H��)��ɉ��4����E��T�Y�p���M�=�஌S�@k�v�'��̮�*�z����\�I�V��{a^��*�j�@qկ�<��U��<7��R��:	��%ȹf�Y����O�JH;p,���[G��r/t�?�Ek�|I	��S��ZSw4��'�{ׁg=��?��J����C��ҀSXO+�k��w��ie������0�u�%����OwW��$�2n�U与�Y�cl��KVU�­�}�����ѪT|�������E�����P�*X�dA�^�禔377ϖ�fX�>�~�L< T	*�!s��VP>.���jJ(��D�h*$ `ٍIj_���3�]��^YWW7w|'��v�B�)͗OF;������t kb�wn 1(-о��j|�����7�ֺ<��F�<�*�dFe2�GC蔊n���o\�(|z���0��L����I��wt�Da(���K���zD�~gC<�e���t�eй��C)%ϔkr;�e��`ֆ�'��O�fFm&E}��/�hg�p���[�<��,�����/$��0�xb����}9g𔨇�b��&�X�kC�r���n}S�ԿDLtai������kj����������RƘ��3�����9���P�}~���uS9Ӝ����h-c�(ط������
d>~���`�u^�6m:}�L�*�Ģ�;��3�����x�᠟��T�=>D_&�����jp�,0b�����ɏW��H$�&�<�/�j�6H?Hes|
qP�eͬsQ<4��9�R��K��;�j�#�����',��ڦO���(�ǎ��6]�k}
����]YYM�U���?6A��р�I��<
�]Fb�,���y�hO�q'����'/n���75����.�b��J�HB�a��8�}ۄFA����w�ϟ���N���9� v�]�1\�X��q�d���o{���|OO�±��S6? XM{��(U�3Ȁzěn÷�|Z� \Tf_��Aa��~��Ã`��Cŧ~���ߓv�2/��K��)�L�{��,!s��Y$�S�	j�1Ϟ�c��5��ꘄ�Ւ�Uߊ% �D�b�H�"}��#��A������� _�w���`ݾ�+�WlV9
#g[�0����O����ir��������s��s�!��0���yE����-C�8 Rn:,:S�
:���ӧO��|�x�1�}Hc�1�.վ �A!!�SChӁ�1��l�`o`0���RWD�ْ�>_,|a�q�=6�,&������D}N�(-qѵtk�|wA�����b��H\���Ш�u�m6��pnb��}�Ԥife�ڽ��G�z��-��t��b���ׯ��Ret$�#0�\�8�1I��z��PaZ�=̡Fό����x�YP@�	*�Z�{���P��|���|�w�ڋ����;�^rs�1/{*fq��u5V�
/b&#�c�=D�>&��2 4��(]p~�+Ȋ���K*k!X�,���A_a#B���޽{��ٽi�o,�Z!�y P�.lV�����d��ƅ����ץK/!��kP�4��-������E{v��$ǭ���t���h��\|��5~v�E�Ԟwj�K��K�����Y�VKHa�
kc�����C��P�/�����s��B�I��M��ÿt�ط*	��s�(���2NY���|r.wg��&Ar���s�IJ:�{���l�z���F�/4��<�y7s���ظ�S�>���TFc���? կ�B+Q
PzCZ$XN+p���_MuZ��`^FNN��Q��b�'��Y�yY��C��\��N�)���>�ym������;�T"ы�K�s��5�5��tp�D�/�X���N�\U���� ��a��@�ކ��[�</�\Tpr�Ԣ٫�F�%)�r" @�&ا@��s��=MMՄ�A�=v�׊���������}�����k�)�i�O�7|rjgq�k��@��R��&oo�̆:�˄�T�7����ƀ��c����]6w��-y���D��=x1|um��P��ġ��xf���	y���3u!���߂�0�z��ΰ��|J�w��4�'�ݕ� ��	��Ί��~2s��lć��
`��ҀI���<�|�_����&���\�|�1�K���)_�hx[��Y�V�*J���>��@��z�Cw[=�F����L��xtߑQ�����߿K s+��c߾��T�(���	n�~d�6��qL̡��x� �p��'�)���+_ZZ�UP��`_�(�$�Ű4��;\��2fyio�}�I	�������c��s�%�>�i޳kh�df�dfEu.8f���57�]G΁���U�1w����y�y�l<S76N,+S�a7ܜ�|h+�9=��x�O�8 FX �
�L��V�b<r�'q��)���>��^�"���� ��8���C'���O�뾸L+���QMh�����'��Sċ9�c1�l /�~����LPLLO@�W�]f�I���t��˗+���r�M3��=Q1l��:l;���` �X�2�A���3�#6��a��T�Wޫए�K�����;��-�o��� Г���p	<s(	UG�=�Ԣ�lܴ|A��u`����Kxf�ˬn)m��'�}��O/ߺm����k\�(�8��14�0`oh^����'��i
�>���z��B���w�p�pN�v�� �m<�>}���ns���#)�X�︊���=W�E�B�qW�Cc���L���N��;��|����lD�ٖ7X{g�	�IO�!1V56&�?��O�1�}������N�$]��r����:2~�������3�z%D?�B^'7:Y�k���� ��'b<��l��S�U#��q����@������EC��!#��C��'ΑU�*��ij�k�4�i=�8���bA��tڿJ�KZ��� ���MSȾ��9�H�RL�b	|����/���ȿf�^zo��]j[_�H�j����½]�q���N�'�2}�i6��c �rǁo�+)IU�׺Qp��3M_�k�y���̰�:v,���M-]ݧ�M�:�[�7:Q��!1�ͽ3� �½vVç�I����G%�����p���_�P>22R&��?��P|�)B82!���df�g�ͧ�Ok�%�~S�����)�|�����f�����>&�|Y[r�������C^������43sjǘm#���ϙƾ��OS��%9
 �⫪c4�����dUWV�_9�'���H�#�e���0':����y=��@IԦ+w���#�Ꜹ�FΛ;�����.~����� �VS]I���W�;S���591zo��7��J,���qjl��*E��9Q3ā�z�P�W��c��pU�L�x�=	嬬��!.$���X`V�����O�� u��)�z�\�#��E�@�1�GkZ�[tlG�, �<Р�M������]��ծ��Ճ�^���4��u�j%��
�z*sC�'����)=|c�!�]�~��%B��|�Y�zW��ĝq��p��[b}���EZ��˵����Wd���*c=cUF��w]�Lg��>~���<���MWel:	�`��S�l���`Π;w,���=q�)a� ������@X(7��#`�a��z����{��5�������t�]߯���+�q�c9�oii���,!1��7�
ֆϝ � ��RO Bifn�=l��x�ڢ�Qh'����6l��̭Ӛ=��G?�
�C
�s�����	Z�l|�������l�j�'0��K�cuM����;�Ұ��_iS4�cJ[��ǋhZ  j�U��d������M�0[q��TEO/75����XS�4��.R�gJ(DOo��������5��I��TjF4 l�ܹ�[��}�����k&-~��$�����I �)0�[�Np�Fn~^��G��_�~[X��\Fo�'y���{ϥ�T���թ���=�\֝��X�u���L��c��/k8Ԙo�$�tܽƉ��7k���ڞѬ�o�! ^�u������V�Q=��*�$����<<^999o��9��HAf);�����ʰ�&�3;pz���6ױ�"��x�.[f�ݯ��?0|l#�y��Ή1
!	��5]qn�iI�5�	��wc:��܆r�������D
��4,hd�5��%s�����l�5k�=z���Pw�	�ԛ�<Pq�5PM��Qs~8��H���&G��k=�V~��%k���Z�*jk�"""pN[8�b*��	��,/��t�p��Ȟ����p�5�uRΑ�$��� �1+L���(��}���W��i���;w.�40&%�R������V���/�x��T-��z4��}��W�h�`l�SO�Q�[j��}r���(GE�%K����⒒ѪBBk݆N�ʹH���AdR� �M�T�x2lm"�C�3�}b�yb�#�ի݊b��10"ҏl>y7ٜ��E��H,O�����~u�Z�5�<��,i)����5x�'�%������/��F«tAL�I��
.y`���-xuC�9����c���'��I�^�Y������z����w��?�c��,`�.�'�3t2{����Qk���p]� <5*㷆�?sVC$�w�^�����8��|����97{vvw{WTT覝�*�'!�XWKT4�L��eR7,=��/�X�f�*�	g��o�Y�8��r���-^-_'~|��tU�����h``��qWM���Fe*!�[*���}$�}j������|���S�gL���;�:B�DqH�_������Bϟ;�������Ñ�ݩ�X�/��_;q4%
S��̛���*���e�r�6���S*��Wnذ;|�������mt�Q%�$�f������[K�^������jM�8؍eY����	���sr�'��=�ÿ$;@%�!���]�}���t��v�n�H	�ft�-��ڧre�{d�Ђ7d(O�(V��Ek��c��ݴ·0�����7���@��������,��P���ɹ= �P�m��[���ÿڎih��.�;;6�!��8oi��tDޕ���]�%G��@؍��<�����*��o�!F�kǚ�����8l�OD���7tfzWӓ��&1w⢸�D��G}||�<�v���&��?9�CNN.�x^���������ud/x��r��&���N��:��t��.j;/��!s��IU8+feY)�-1�a�xkME}�j��Qѥ�{O�˭�wk���+g�\��O�t['�]����F���J���h�0���?_�U�] _
a�lr������v���G]Z���/�ǃt����m��&ɐ�����͠Q�
rs��<�P<]L���U��}h�|F��P
�+Dn�/�j�-�"?��(�����vq"w�;Rޱ�"����'Ё�}�~�Fy�OmY(��j��lrc����������I�u;��
�	G�
��FIػ�߾��V+Ry�!�j@=5=�]���]�V��<�!��D��HEc-K�m,s�0��fů�i��8�
&��߉��:���������ٺ�Ŵ��-�E���ƙ������W��d�+���8�_4m���<Ϙ�N�M�s����':��V�7��xr����C?�����y/8�o������Ԣ����@�bd'0�M���w�ΰ/^\���[�F�1tL{`�<	�C�-�`�R�'s~�#�������g��Ƿ�>79�[�;�>�Ym�R��%rw�[�~�N2R_�T�E���g�5���|IFfr L����^J�p�tG<����|�3�9:�}���u��Z���u�GF�ۀ�D/��| ��z�*��8�������|��h�&�D#�I��6���f�)��I���</�.�lE(-Zsi�v�!���iEc���{���@���� ���_o��^�y���+�d����r�W'ˆ�Z�[�b4b�� e�ޏWz9���HL���9�}Yפ{Wk�ހ"�Ы_oI�#����d�N��)��#$_[�Z�U?��i��1��,������ϯR��?���C-̟.m���%����x��s�T#fy4����kݸ���ϡ��bA����ɿ��&���֎T�C�n`�x�LQ�|= iM�?����/}n� �* �,������osfR�qп�5��Sq�I�GFG[�B�U�,K��q��	��L���L�Rt�<��0��.���J�po�QX�R}m��,D��L97��Q���|v�?6d2J� ��X=�r���d��5�t4��3�V�!h��X�SP�a!6���6�"Lf\B�.���n� ]|cq���o5���0
�iu����?�����A��<ΒK�½��	���\��+3!u�7����^0�-����s��A���߸��K��<�MYD=��@9�ļ>dz�3J�G�풓#1l.X~�p�p�~+�O�nW7�V���iI�2�	����$1+�WO���:3���-ɉ��ʐ�Ŭ (;[f$ɰ�gӯ¯�gct��5�t�̙�`Bc%�S��%��IXkc�>R��wf ��i�Mˣ���	��3-������6�d#��m�xӔ8�e���;,8�fz�.
�м2��9Mgr�^��n{�Gm�����?#k>�O�:X�ŻThsٌ�44-&TN5���?��孃@~pG��.���NL�����1�Y�qM~�m!��٘�ɷ�'��j���8�r:�X��N��-�m�8�6$te��*8�c��FAo�m����� ��0�6�XAw �?�?��؉���&�R�=�>h�cin�8	���>TU������9��C�2JvLq�t�m�BB��?���.���.�E�S������G�SI�0�L��o�1�?ZH엚^~P
�<���@�UZj*�@h�~��S�J.f"�^��Mw��N��5�����޸v�Z�?��@�o�8�5�8]�
@�N��2m.�Q�G��ZM�*�9%A��\ܐ�}d�1k���3�Xڡ�>(�R8[���%�	�u����V���:{�0�>�i~��a�;͙���������刍߶MM��@>�5H݂ �.t�"�����GsY �p�C.Ғ��t�^�M<�-�^�5.)����JD�"���|��
�[��L�3�m۫�*#�N6�	{'2==��^��2ߓIwILe7������y���`Fƴ�H��2*8:p�cF���Q�u�uLBB�Lt{o��8��F�X,�<s�L���bH�+*������~�.,X���}���OH��RQ ��U�s��)%��|�4E\�oC#Qm�k�;%�!օ����7�2�K�Ȉ.��6oR�M��8���Be J��dN}�FH<U������v[<}���^VB+��K��n��=߿�`�M�
�<��8�룋�ݳ�KXe���������*�Q��8u���kl����_/!V�yoA80*z�5�ʖKz��Y�g� q�hR=�����=�{cc��NvO�.�P��D�mZ�~�z��23�a�_�P�}�_2;����|�j7�#{&?d�>aaa�1�n���i�ijr-�8���!��;χ�ڐ��`�z��0Z�2A4���wV"Ȯ&N/����jz�$�
�L��&�M���眜������{bFL+�w�}���I��ro1(x���>�`��Q}��tEC���]�`dF�$(I�7�fJ�*Fjjj0�mF�R��*���zW�&4w%N7Tlkj
Q��Y�^���u}Dq�[���g9tDMk�-udd���ɽ��Aڂ'@+�b�t�F����ψ�l������қ\"�Tl�tT,�6�|�hu6Ǐ���; �@e�_��L���0X��zw�h��<�����+���M���c���] "�q�_H�de]ݪ���(�uK�O���.H9x�!��+�ٶz�� �F�������߿�  *FFn������ G��r����͞�?���l0+k٠B��X:-S�T��"|����D�=|�s�/v.;m.4���i8Ԉ�ݦhllL�hV�0���U����*�]ӟ*Z�Hջw�>�p9�������'����ʜ���b���9=0� @xA�ϟ� 5앥��sgZ�O����Q��d�{�R�VΛa$V��W���[b%�hق��B�W��9���iS�t�t�fP0õ'�"�;��A��z("��P�THj����7-`�T�ȝ�����-�M����߮�6w����/�K��8)1?&�˯US�<���\L��.�8�笀�r��g���}o�Vx�����!u�~�����L&�s!������h[�\�rl�Գ)0T	1{| ��>�aqέ��K����D���c���V}����!�!e���`�LN�.����w�]eZM��[j_�|���� ��@��ݻ�-]j�ċ��%o􊔼�n෯W==-{n{�L������*������/o����h C�TZ	tٴHX��J!��Ȣ�(d	�BNjZ�'''�6�웓�cim����677�ئ|�ĵ��7�OFc�>�Y�����8�t�>��D��<�Yjz�N���ģ�`�[!�E�K���>x��V����������@20��@�f��6��py^n��	���^��0�ǃ+0:\��o,\��ld�������t��.2�,-J"�#1�_��Ѳ���B�Y�ظ!zC�Y�B&���i��u�G%�\bH ?I.ÿp�̫%m��O}rA�qn�q��dkkH���00�6K:��_XЊ\~��[����n�;@Б`������o@+��s��n�A���&e�/����V��#���zմ���@}l'��K2ՀM��T�]h���O�N���d�v�a�" 
>�� <�M��]]^���0��ջl>5q.�r��-��-"B�q7����P#`����]�adOOߗ�S�&4�X�D?�����|M����>}�E�_FP��B�l8<�s���u ;��e�>q[�&����x�A=��"��í��o��ˡ�r�\Ļ|�s�mK���F0P�B��������bw�������mWˮ��7f?D�gF`X��*`��l�Rg���:x�D!�� nr��6�7�[�~���g����-y<�a3[0��n��>���Ba'k��e 	�.��\	����I c8���L��<g�i�b���zj2��́���2A�b�o��6NhR�޵?FDX̝��4-��)�MgO�?o�Ic���7���_��Jy����jժ�66��R�2N���v9�PyT"a.��k����\�����&�
�B�T2;�S���I�<ώS�Dʔ��$���n��3�e��3�w���������/g��s�^�Z�u?���¸�vsV��0]�jK�=�qp�p!�9�����\��$r����� ( a�{Q^��"�9J`Zg�WM1�UeeM
v��ia�Imu�A�� `�/
�X̢-�*�C9R2�>�2ӚW�-��r`3sss8��o�'���]B4Cv�^^�d
8~��OY�cT�)���y/� ����h��oݷ�>y�d/Á����J��-��X���MB�~�ԃ!����u�Rʏ�J[�d��OP����)���6�*�i:���|^�Ao�|�c�Y���ӎW�<�ry�-e�Hi	�ŔNH*6t��;���A I��>\�'��Lu�&�@^���-�����wu�u�I�a#W@-��34�wY�ms-.�6�nhbT�jaT!w�3�1�,IZJǡG��:�Z�v�a�Q��k;�I*�O#S�Xhw% ���4�CSwc�Xx�i��x(\���Ҳ�j��ȹ^1���
�5,,����w@�9���1�8�%!!KΥ��j�Fr
-q�%�����!�:�_�F�W��)Sdɢo�9�������e�e�s	|��W��k����,�� ��̀	d�$t}��5��]Gk�����D�x���|Ȉ#w+�'�!++�OmP��ò�%����16�\�Wu����R���S9����0��Z;(����y|ͪfa�Yp#���\˹~�$ƗqdM:zzy�ڄ��WS����7cjkϓ��Xr��� 3u����G}�Ʈ�Q��x��ִ�tͅ��=����l���~�@�Lk1U|����GC� <��.-=�e˂���?e``��(ר���]�lvB6ݼߕ�M����rճD�q��jvߑ��!�7��(��T������ݳ8+I����	qꍖ={�����ft���*�qqq�x1$���8��r��EY��+��`{��:�:�q��&^Im������7���-.,���@+z��������t�+[�J�$��a���'wRT�BU�x�:.·w�&�S>�Ҥ�˷��kt�Y��N1㗅�/*�����K���9�g�����\c��Q�eEL�����M�g/0L�#I @�B��!j�OIr�Ww�������M���N��^
�#����h������I7�/��|r��w�L�<A�*~~
�YB^�͐��/G]�6�^�b�l7��ހ��&k/��Vn���b�uh\m0��4D)eO����[��&o�hyww���Rn4e�UW��xU���x�w��ˑ�%!E�G�� 0�`h��Z��XA�A�".�N�Yʓ��k8�tB���餴�a�s/眡9 ^0~��w�_�6��3F7+S���zr?�)���⓾�l�<A\��ek��g��Ţ�����Fm�]��0V���+����ԥ�5������gl3����HW��;7��9�). ���/�E|�);�f��#WUU�_Us�^���H�E�i=�n޺�T�IyM�r�����[�eg3::�����I�㫸!��%ෟ�(���"\���P�,���bZcT'�Ny� 0�8����7����O����Ʌ�,5�(���!`��ٳȶ����&*	R���ױu66�=��q���%�]�aE��a ��7�Nn�~��l��^p�]滇�b\��R��Fݥa���m��\w'���$/�} /�H�1ta���ج�f��O^l�5�|�^l�YS�\ t����@�cR;�Aoˠ��T�:ʚ�1O����--O,�����q�C����ݔ�S����SP����"q����a����~�F����TUV�ƒ��o� [��i�[@Bnpὥ�]��2�����X&Ld)S����,��/�5jи�+���Sa��--���\��qǉh!?���C�D��C�Qv�r��7��{M�[����7����.��s�n�̱jԨh��?���Aު�7t��3&���w�#� P蔶G"��@� �a�v\����_�(��"ۦ��>7g��аPW`�U-�`�]ܖ�R��"OKؽ�yX�.���L�w��z�|���o)F������5��-5�EFզ?qq�f���<1������ |b&����GiC���W q���
q������Y:�~?nk���hB�235���4�EȺ����0.��o���`@�}��$��quu��y� u�d�P0lѩ���'�1;�*r{�ې��w{z»x6��J8�����B����(TmC�	+$���I�ס����� 5�a^o@4z������5333����yy�p�3�zAƅ����d͏?��&���O��3�Z�G�[�Y��k\�-��Zs�Z�N���,)'k�b�Rz�毄�dPu��ٓ�
�8�"bA��$��	�>�%��i'CC��C��ۉ��� �DA�^�elll�+4΢}���' xV]A��j$���b��)u��-4#
�%���^s���U���*�5�E�j�7��fh;#�Τ۵ ю�)��m�=K^���-�h،����(�j�}����-�B���k�T�\�y���^�~�ݘ�m�O��!���2V��G�#�����W�I�M�B�d�+��E�p�M�.���^W�3~��n��D��dj���?:
M�Țȼ��Pʰ4j���_^.C�ۈpxP5�(� ��f�f;��.�d��SVV-=�	>� �H�@��W�7��D��:�4;9�6�󤘘�<"֢�Z�#�"{�����	���f�\�HY!I����������y� �,dl��
�@7i/-�,W���?&��pp�Ɓ([ �-;�w���d烇X�`�e}����P.�6�$�����.BJ�CI��@࿦"�-$GV���5*K���͚l��ic��_8;5��D�~��D!�=kћr���O�Nۑ"\�����7�����GmB�w�G���P�^��*�(��,۷C��GE[$	,��i���Ve� 	0j;�r������5���``N�0� ႁ�<�Z����D�N�iB�p�%�R�^;;�Hy�[��'7�SfV�҇�yڨ�*!UNQ�y�Ĭ�3hܳ�ewvv�@�nyz�y��/�y, Yʏ�t��n��
�����@\^C�Ӌu?pB���ID!;����܍������b�h�3;�l},�����F��Ƃ�'����(����BhZD��A���D��ᖁ����^��A�w7��mも8GCk�Z�g�q�^PXD����Ӣ��,v�����G�!Qÿ�t+�zv �sݸ^BRtS��.B�H\��+�L8s��a%W)��I!O�0����$ ����=Z�E�u>���9ȢI�aq_lEhl,�e���l02)�}.쯿�"�\yBE���3�H��ʲ>n�0�a^(�ښ�h�̶�R<�1�v*�.�#E`�
�9'׋1Q�p� Ty+����Y���Ť?�Mc|��ڊs�Д�ɔ�ag!�S Ehs��� �	�����ؼ9"*�S������CD����m&�g��Ͱnjg�^����6���yӄ���ڹ�&]%}��O�HJP��W�������:��[��]�*��p�^��a��B��U��'=�k�^^KVڹz�L��>N�s�R�:$3-qf�a����ؚ����
l8��t��$�~�4n&x�̸����������;�HJn�d�����_�˫��O���653�DK��B�	y��͛n�PfoμW�1�d]�L�{������U�zzhi�b���|cpA��7�O-1 ���/υ�7~eQ�KJ�L��A.x/p*ـ��o�k:fAL�'�����d>az���_��
p�4&�L����׍�࠱��.��S]�A��J^6��P�]��4����~���YBY���˗!{B������A0�|k�<��Md��틻�!�i��	a2�[�����K��K��j�s�!�F�3yS�@�[:��y��9{ԯ��Bl��7멐�l3�B��_�>ыI��W[�j҅�F������,6���4i֕�oa�e�s��Z�����օ����ߵ^|RS��E��8�o=�ɵ�&�lVW_�%�SJ�����%�CVRJ�3�.a�j ����)�������	�� eO	����.[L�S,B�Z�9��>݃,�5����ӳ�F�lS�9�/����ޛ
�k`p����t��i�	~|�ۓ���(�J
/[Ԛ����P �<� �ŁB�DO9�U��׃«�Yy�{v�G�r?�K�ý!>��� [t�|���( �-"##�{�F�a�h/*a��Gi77�pj�o�/����Cv���>����������;����S�����k��D�����`��e�4x�y!��3�����Pг�v�_��D|$rr����4�ir�HS������;uOI$��'��č{N��g��v-ҷ�
���fgvJ�l��f;�t�G{�ns[y�:l��+�&�~Z���~�:�����ނ:��إ��D��"�wڜ\AcM�VT���o�� {tK�?ioH5$�p�����{K#�&�X�������fo 6�Á!�9�����t7���W=��+"�^�����p�1�����	e�[`�~!�5�߸'�vm�a��;Ӈ��Nn��#e͐�\ٺt�֨����_B�ۏ�>ccc���{���W���b�#AP9|����4�?����٥Pg��)�d s�g�"���v�>��M�o|�����/>>�v�"�8B|�Kym��*K
�j�)~�;L$�<:0e�󬰰���x{U1.,`^)&�����1�>Pboo�-y$������Ե� ��<���(���s~� tZ]�ABF�C_����O}d��,{!�\6�����!�]�^f5j�,:�������H0��"�wKE�,��wo=G0�����F�[��+/>F~9?B�PPP`�i��0�֭�?at6&&��޽{��D�� ���؃��F����|��w�D�����S�4���4s;��g�����_dU�:�1Vp����D�3r�/E>U6�<6ߪ>�!��a'�+�U���T�&� ����Y@@Ey9��0�|����� ?Sè�)�b�}2�6�"�o�q�b�~� ^Qm\q^0\������n�=��p����T�5MM����A����<<&�l�^[[�Lh	�o{wP9�`WIH	�`n��f��x?ga�`l7��c�!��+(��R�A<���Fq�Q�`pk���OL�n��r�x���uȫxf�جg�O֪�qH���l"IP!�ߐ��,�~�T'vAgvrH)^Kz��ا��HY\��Kb~
R�����O5��^B`����=�|)b��è�T������&�4?
���%,H����/E�����)y2+����x����D,u�3@^M�L^�0�=R�
�;
L���'���oH��Q�o�q�@�sI0�����n��r��&�	��@�0Q���4Y������xw��9�/R>b���3��_<�=��HoTl'�N[x9u�<#p������>Aj�N��_�S@��W���v���<�����D�^��
�1�_b�?���$텪�Rg��b�� ����!��=>�UңL�LO�Q���_6XEk3�J�V�����&&&�����oU��cV-N��cU�?�a0\�Gyno&�!o���czv˝�A4Z`s�Y��旇�ώE}ݯ�F'N?��K,�%I����Z�C?�qx��R6npݕO�F�W����?jѼ�
��8��e` ʄ�;�~$�dAU`���l��>�,P%м������׽W�S#�$���H[����羢@���|N`���`CJ��y������U��V��U�t[��y�c�pT�Ƥ��D,��غ�С$��Eqd �Ԗ�D\��޺�)��v�lllf��D��6��a�����VC�嫄K���v��X���3�Px�Y,H� �U��⩥3�@�i��"Yd i@D1���G��w =s��
ѣ{�]�jR?�J@r�]�Kl�U}��m(b�s|��XlG_p���駿Y��5�l��]�3���oZ��'�4:�@y�Pk�<��i=֓��xwŧq�����%�JĎ�Y��X��G���3�r��J��.��/ y��B2>Q���v���p
���:��S�_lH�οU�&��N��fVo`���n�ϫW�p},$|�tSiIUMM�Z�ɿ�����.]4
�.�;���+P�!L�A���B�C>"���R��h��q�P'�}[�	MR����Y�� ���>x)�Č��At��Kn!�q������5�G@����p|ρ\C�1����,���;�531�0C����p�0��fL)�8'%%e>Ф
=Z��#�^� �	�g-��T.�{�����d-�D�"�2 �lOY��"�0v�������d��h�]�iRn�9��k��\�&L�y�?���f
�\����ʪ���Uʹm�v����vN�<yY1oJ�v����-T�h�VJ��%h��ޞ�޴A�c"2��%7�+���ӊ����ۯ�=	�6)d��c��&��"�B�����#�T��ROT40�222����/{;˒��gjKn4�A���|�͠�M�Z�jk�qE�G���� 0��=y��jbLMM��^/���1�|6����!~RA��xG��Dnh
��(�@x�TZVSS2���[}rW����aFډ� �%�l^{�6EPI�F�'�H~؉�PJL���o�h���|�8	����sD�,� i�6gcc�)���P$�P��I�yMڹj�̧����|�f^J?9�sE9A���`�@O����o�>��yyx�b��b�7���m۶�o���f&��&p�U����O�O�4�)�@�����d3!�@@����4�t!��jT}���p6�
�Q���$
��OdC�F�`�e� �>?9"��)���
�7�yTP+ ��V����n} �G��Bŭ�1=Y֙`]����.,l�Y#h��s�QMooo�Tcmԥ�Lđ�6�al�Yq)�� �`^�P�?FR����^?�PZQ�Ѷ���}�.�rU�!S�o�,��|
dW}�em�����q��H����ʤ��V���
��y�" c�p������3\[b<d�2�A�ݾ�8M)����>���K25���-�+��,�;��؅����T�8cc�;?����~q8��\�x���Sȴ[�LZr=JB��.tv��ܔ�}���E|�S��H����f�ׅTVW����Z��[�6i!���ë��p�B��.���鯯/���j=z�����R6�w��Hun���\�=��X�
V�폌�.p�6�b��R���c��7LSi��	�dJ�Y�|�/>]��p���SD$ip�W��I=ڑ7Ԗ�vao9��q��dd8�1<<<�QRb��c�Dtt43y�Sٜ�;/d��9�@E"6f <���s��m�st��O�w�����	2��V.���� K�mO�7�56k��<����W��!Q\�E������L�w��	�����#�.�h�b��8�!>�'ۉ�Ɨ��n�����3 Ԏ� �@� g1s��\�>�>?�=/�n��-�z��'s�w��&]����R�I� Q{w:��@@b�X����i�jbe�tK𚇡֜�o��><��K�C�-89q>�x�c)v�������<�O��o(�H2�*B�:��hW�JG"z
�rqad˯���
��8��g����$�FGl8�h��R�$�F����y��ā<r�!�0 ?x�j�z a�o����@��c��F�<��OVS�#�%Z#�EPK�\L�t/V�����#���ő}�3�qf����C"O �	����5 �WJ�u�J���D@I���t�D��a��y�S�Ne{Ǿ��!нʴ���)�K�I��G9zo��W�-<�]�/yK7��{֋�)	>~vWȤ����Uk/q{77u�JjL�r w�L�06<i�@�Q.��K�Uf�_�t���+'��Sa8�e�\⃮z�]D��g5^�3�y�l��8�S]DǑN�6�t�@����^�k0c�3�i��#^������O��N4�X�R�f7��@��Px���VEA\#"�{lԧ -hP�UsM��l��mhr,p}���,��=�>�N���'9��(��$dV�ӫn�aV?��_װ��v�7�.4/$�����	�~R3~mV��UĎ��ԨUG���d�2ż��>,=]D���en���92�4�GP�����mO�۷?�E?ĂlSN�/zvLo�O}^S�zH-��8G�����Y4����q��.+6�0�_�h���
@���c���H�A�Y��!6���"��HM��&�~"�s
�� -j3�LԬ{�q˻����Ǯ�@�0\�Ϡ�����!ߛ'h�QAA���*�d� �F�#8+�y)���NN�o���� �I7h���Xz��V�Aќ���fͅ'}\�zյX��& �Z^�/vٺ
R�e��\����`�NT��zl;|�o�	��t����K'�7�S7
��ޜq��0�/���i2@لX�*� `c~S�M0(�K���x9`i��
`,��X�\]�>��Ԯ�����m@"}��F�JJ@
8�gq�1h%��?�(�ع"��i'�ֳ]�!�?�W;��%h���^t`� ��1�],�����qJ	r�����H�>_� ��<t���_��͋( '���y��=W�����!�m)�y!�y!Z@K���9���g�l�
�C�I�5j#F�9��q!pK����f�t�sF,PK<����]f��yr2s�Jf�U~����m�S�L��o�+j�=���d��ma�	��ܞB��B����z��^�%]PP��usyMӎ�%����vf��APǖ��s�|߂�C��x��=��t@O��:�kY��)L�0�x	���o�fpQ�����}.k�U���D(pg�THB�'4�T��-����� �q��6�w����)-V^�W"��|�1������x/C��	r4`�����^�\�wI̺���von�<���6"�	��ː^@f�N��`p�bQQ�UbM�f�#<W��,oNw����s�AF(~��p	��ϑ����;u�N��^�u% U#�|:]�A��m��!0'=~�U\\�5g�^�10��� O�k����P�^���1ș~�H���X4���Z��5۹n�*Uh��Y�e�c^�QJ���{��RǪ�M��F���WG+WTW_1e��I�������q+R5%�I�s�Y%V#ͅ��K���Grc���ZGr(@'2/�Б:�X\�[�����M���8�%DN� ������9��O�AD�W�*�j��vs�XWI���=ni2�,���������|��a�@䍍�����L\���<��J8�= �:r��@��?������3����1����z�������,[^GF�M��.��5�G��������v�k1�C/]���ZgkApiiF�����W�g$�<�K��8�E��X��\�t�~�Q��):0�8��'��H�~��#�]vX�S6�����\����/���逵��b�&^�sL���2��!4�cѢ'�h;0�^]����x�I2�cйZ�o��O�S�Ĭv��!V���m	�}0�g�����^�*�@f�A)"�~����X�6]]]��w��M:ρ6Y3)bi~��.�[�wcmt����E4@���qڝ[x��:!�NaA���_�*���3j�g]���r�*�a{���I%1s� �\~GL��c2�)� @��-5ʻH`P�qd�� 낂���E�L��}��W		𿙳�c9�UA/B����3຀`������A�+Wn��DFF�^VUm�?��	��U%%�����i���^ 
1Ԧ[܍�ٞ��@� �Ԭ������g���:ǂw�Y1����6y� ��5����]#x�~��A	��K-���P��t]}��t_�Ns��ρ�|�JV�0�D�����@�O������6��M�J�DP7��'�B�k�Q����Q��H �_�Q1�@GVU�;�ׁD���:	'�\�G�(�^�O9�~��D<	j^�|đ[�����j#0���U����ٌ�P�!0������eho�eHp���y�j����~C�Z�q�� @s /�7�.s�'k�kHOK����~{5��X�g?	�`�4~�� ,�']�l��q!(m��~꺪��g���<�����ׯϜ?_t7Z���
z7�Cڸ���d4멯/s���d��4k��	�֣˷;8������<�Ĳ��g>vg�;�:��a���2�.�=����#�˗3;��E�/\�|���
'� ��w&�QVq۔�j����Z����S�tQ�N���׎��y�3h�@\���d���v4�˃�n�]�߆�?s��Z��g�(��*��?��ϐ���7�oKA� ��Ѿ���#8�0~|Sf7[���,�~o���w,m�QCY��(E��g�����FG`J[c��4v�1m�5+U)tN(��|��֋�ڛ��P�����ձ���*'��h�<�Y�G��/�ߔ)�(�G��Wb�{����3�j�Ӵ�YRt$�aЗ���T5�h�$[�^�}���7�f�TY�eo#8�h��%.�K�t�9ٴR�1��x����z���9�a/��GM��3�9�؊���+�8�V/?#)Q�9"�S���D"��X~�t}���q<�C%*������(�f:������MOOo����6��/�T��JKKn";�m�Z�����3�t���~�J4n\�X>�	�!7���p�r��$.�L��u�k ]�VwP=p�'
!�������H�:9>�w=U���G�l|�I;�oY�&�^;�����ˍ���� ^��i�v���7��`0�l�XT��!@XD�f�8�m�0�Mu�x�ML�@uZ���Z��C8�Șiܯ���3jB��TM���b�V��I;�,�ö����L��c��uc3Z��%@�C�TL�
�P�Ĥ��<ΐU6��ĹҰ�H��{͗�!���\��љ���S8��r怣�Y�P=$
��7{V;�9B������ t����C��s=��~��&z*�l�p	�#��'Xv����^���'6cS�9@�Lk3���9V����<$&�n7Z&>�}��.B�0��W":r.�1���F��"՘;�FˤLȳS���h'�NՖ����>ק~��:#7��8�Y�|�#��؏'��S�C��n�3u�AYV�C�&��v/�N L���뛙ͺ��PjÅ���W�&�@"�O~��j<�~��s�)#����!/<7�6�@}��-����� �M� ��Y]W�,d���nc�:C��@s #s5�����M�M0�	ҳg�Q�PW����ꍌXs�[�v��L����e�3�������"�`����ٿ�ĥ���|�^KSU�7N�Z���5((�)����?�0��moWF��'?b������%��$n�q+�z����C<P���e�õ�����}��F�~)��
$<5�ŋ�O�91�+�jA ��~�Ձ��"�l���\���:d���Zl`/�����/������޳����@�+����\��`1�_�̄�pc}5�AC��爙�m���6���i��/cx��is�j}��ky���)	!�a-x�$ԋ��k>�z��%j��ުS:4�pB%k�� "!!aiuei:~�&LEeOG�ZX0��� ���_��@�<yb���G����!��&b��awf���X���܊S��S�b��KR��)� T�x"���dTF� �>b{�M����֡ͽ$R�E�H�k�q];<
$�	��e�/i��X�=�kq�^Zs�����_�3�-f3���m^뺝l ;@�/���~���w��xrvD�sy�ZG�;�&&& ![�{]ʇ�К1�	+�~�fD̘���藪�$����\�)��?��Q��5(j�K�!�n�i�p-���ˁ��ƥ�S#]n�S�<~��͎�v��
��¸����s�b����9}r����_#o��YV��/�=� @��b�K1��4Ϩ����aI2�.�ʄL���~�.p��9nj`~.���_`Y�`���^�a.v��YX޺0td�)�1\7N�	�~�5����0eO+Ld7{i�z�+�;�4.��"�e\T�ub�o��������)�=�ů��E���`�����9����p�}��@�sy�'�=���;]$f���f�(��|��)��T�
�_��m�#�v<�ي���aX���O�P&T�,?M�g��.8�n`�?{D���cf?��.��y��Pw���_�S�-���U�C�<��M3��؁��o&�S��l�\�������|��� 
P&�R�@���`xv��9�L�^�j��4��kl���X��'��tEFs��]W�dv#�ƒ�E����C�q
�>$��������y��.�[���s/�zJ����w?|	i�ܶ�G=T�/�~/hQG@��ʂG�ϞH�l����?
� uCX�C@>�����H8����mm�w~X���Q�	��o���f,G�փ�����8ÁgS��뮀�Re��!wʤ*U���U�d�'�~����q���(�<���7����g�j�[�N����NX��
�}�����t���z�M�6nz�f�|��2�x<�!�EKϨ���]\�ݵ����j�5\d`/@���Æ���A7Qkk3fPq6�f�C}�ϡ��B�/C�G��:����H�����yj>�\�������
�f��C�,qf���P=N�^)?��@1SPy,k����i��CJ)��:]�	�}��%I�aLS�nZyU2�^c��k�/���}��������J�P���t�_�{���\mv�]���K�rgY����(��R��H{X|g��2�N�K@jXW���XI�	n,�n��������zf_>u^�}bN3�G����J�����20���O��l!����ƃt7ˊntww���xƐ3���{..2���V������^��W~i��1*�����?~\.c�ӌ����}<�8H�Edd����w:�1�}��ܾ��#�bﱟ��EB� n��%�bTC|��Ѣ�}nf"��]��+��8'������fև�K���U�pch$d^�UD�>q%i"���P�����}��pHto��C��\�/�鯫n�w�Z11��JTN�|�uc�#u��/.E>��ˢ�����a�!p4��#�4p8�e��l3�Ɍ',LOO{�S��ٗ�\�y�\f���]��x�Uz��+t�z����)1j��Цd2�\���i��v cπ�w�Y��"�J����
7�М.hλ����|���DϖP�����������#��� 0`�'+I�?����1?���nsQ�l�[�W3��y� ��߸q�l��#}�$(ˎqMʶm���R�������Y�mR�vp�ioN���}9����ǫW�~����p�8��ˡ�=\#�3����Ƈ����Kԓ����2ǉ��:ũ�N��}�xN�ߜ�V�l�q6��5��Ά�U���]$>8�����s��mLa6e������ 
�����)�۳g����c�aX�9٬pvv�3�)�mk㵩����{�Q&-���LK�g�ka�3 δ��R#��BT��T�o�b���4���@��-�_�1E�g����w-��;��9jZ�N�F��e>l�b�?�Vw���f}�9 ��=�Q��3ý���Y��+&^��F'7���|K��\	���Z>ˠ�*άn{�����CY�ǻk�|�o��2���R�_B����E`t���w������]�O� ���]�d��+�W�pZ�3�I���#d�������W�0� �^��ō
�z£3���b�������K��0�[��w���}�����W��:��7���8�5#�3�n���GO8e�X�ۍiǶ�P���#'N�H�ԖPn� =����0$����o���Ϝ��>�#���\%�"�<���T��׊	%�7�������T�UWo-**
_��� �1333�a����Qn2��GC����X)�;w�|��EԶ�<�^����ge�����b��<����<��ێ�'QWF�5뭌�̓�߄GEFU���V7t���1����a�UR�Qז��͎'���b?,$�d�8�hǈ' =~���[��5�J1�)?R��,@�+�"�UMS�ה:�Gj�O�x��|�n��x�i"�O��b����n2?�=,*�b�f�}�]0�3���f�r*�Ң�30��LO.�����������:�t��OF�=����8���s[�v�/8?_] ��ҙ�hl�<#Z]YɄŵ�
iii�x��� ����?�)f}Wz�D�^a�*2uNtn�b蛦�w�20E�DU�N����-x�Nî�����N�lV�b����啨S��qP$�r�gZ�������� ��/��il��n2:1��׊�>��[{"BA8���l<l�aVVV����[���Ш�����y����	�A�@1��Q�M�RF� ��J�6<_�zv5����	��E���~� ��@��P[�,(8	�U��	���Err��N��i��R0w������ˊmQ���|�ÿ��u���se��©ٍUY��MȔ\�j�,2q��z������O�C=��m'g;��K����]Ij��S<9]��Σs�*:�h��/��H]��N��v�P���ÍKH����R'����9�Jo�8a֫Py+����J�(^R?��g��Km���=D]��i�wK�����=��BMx�iݺuq��'�}�w,$��2>*{|�o�n*+��y!𾿿?��^3�>�t�F��N����t�q���K��oH��ܸ\�0@�Qg�?��E�盪[=҅{VX\�'��)[�I�[c����r����]�^?4T�l���-����>��L�Х��c��:��J�ˤ[Uo�z���w&�rܘ۾�i��ֲB��"JlL�������t��GT�z�.`!���x��I�m�9�wRn�ō��QWN�����L�޽y��A*����q�n��VT��C�\h��f�!b��'��!r�"mGݨ��7;��3�:ϯF��
��d�a,�$PĂ�{�F�7�O�RMt���渭�[F��y��VP~xf�	 ��{St�u.�ݼy���z��v<)p��QZnE�7� ����A;�����eJ�=z0%���8�����������cc=���9�Y~��]��@�����{w��IWq�ؖ���y����H>�	��	���ު(̊W����Xu�u��?oK�@�Jʚ�9 �w0���W��ek(�}㼼�Zx�3�s�n���_ܷ��w����ϟ�X�K�������U�`a�S{H&�''|�_I<|H=K��իxH�E	���Snge�%��g�]���R�;���K�Q˴N=z&*l��w����׵��B����f;5�O�x^0��]ӫ����oRX~lY
���p��Q��'Oᰜ�@~c���G�wv ��9k�D��@�>	�K#<4�A�C@���-<��q(R֎�#NM����2J�����fx�4�-�Hr�����S.��T3Ѯ�y���K�>�zeB�&�g"��0�	lO�=z��)MM̓J��$������^�O��o����2aݺ�1��?[��Uu����C�%P���p�����G�3�B1e�?0�a^^� 0����o=�J�Zu��ƻ��H=Dp[խ1�6���\\����}i��J�g~܃?�p���s�#�2g=Z���� ,�q��@����BɒkVPٽ�!�J%z�K����ȴ�
{/wR飝���?����w����]��*W����U���w����]��V�8_�V�����A����׎$�OLW����ΩǤ��4�+�61P��������$�_j��K_��@�ܕ��-ZMG������w��+�]���
y���!\����+�]��
W�������w��?Vh���@zL_����=a��pqպ�߈"��M�-��IwB~�����G�p�o]߉�)}���1i��� PK   C��X�y�H$  �G  /   images/81d9366d-a3a2-4692-b3d3-374cda370674.png�{wXSY�/$�P4"�A"��	!��� %*HJ��(����FzP�Ti�A���@ $t��$03�{�{����������}�ڿ���k�}�bq�4�g������MO��@�""�Ob�ȵ�~��'߃6""�f����-c�ȯ��'��v��z��%g���K���!����<6?:�Y����ς�-H~s	Q��:�Ӱ�Z��Ml�*�Ft�ȝفC]sGqU"b��Rd��W�G��]�5^�-Ag�T��VGF(	}��Z��P(
��(?�P��/���N������}"}_�A]J0�M�B�77�ͫ[4�Sv��Q
�l��u��STXMM��p�n�8����VżS�ẗ́� �������7�pү�4㏫���K�R���+' �����p縊l���ySŬU�{f�:�$�2�����\ӏ/C-y.[Р��꫘w��!�n�p0BI4�&Pr-E�Ő�VF��榭��E;� �H�d���R��j!��yo������I2�-B��9nZ�\^l�+�l��b�U���k�]���JQ�9�;����$�K!��DiT;x���/�)�d�N�ص�>�e�	��z����ʁ�E��|U��tӅG�����Z�`:��ڭ>�͗F ��B7��!��%��T�6U�ǵ8T$�'R �5m�g�����W��NhV]��&��5�é<�-U��2�xU�������0HY�k!��B�
ل8��o����C	+1�pܒ�A�bH�WC�5L�hM���]qU����
�aU$�6����������IwJkF�[QcW>��7�.d7l�0�1�I�Y��8~��= H�������[Up�$�������A�8ܔ�\�a��Z���W
�8��(���? @��������? @��������? @���������p��ˑ՛��!��!�L��DK��ɿ�K������HHAV.9vOTI�cƻ䥞�"M���Q���G#!�x��@�nϋ���]�M_6����]U�]Ͽw{���8�b�O/�
�1�PF����q3�_:�ª��DH�~0��g�/��Σo��9侩s�Z8�c��	L-���=̃"��%���{�V6��Y����t��ٷ"I�7��%���_��pBklG���5Wd���R�EX�W!H�^�	���Gk�#ͣ(.�±6ho,�[Ej���o���X���#+oK�����P��\ �jC4Lh�y��琉��k�Hɮ@>�"��z���D��Ņd�E;�e%�V�i�X�0!w�?I��"��^>p�S��y}�0���©n�y�Rq�@�
���QT����z�'�b]�Q��{�A'~I�cBىm�W�o�w~�7�-^�~��̽��JH\ :��y&�@���;�v#m��?AY		�h�($R����mp�����ׅ�����p������"�X㚶������F��������	�݂�`ˌ�z��4?�UmfB��-%�l�K��j{͍��G��^u�eO��k=r��\��f�E�p�#L����K���<�A��6f �:)�k���hkK��{R�6��!��g�x����8��E8 Vki4}���4��mØ�����>���Ur�.��oBǚ)i�NX;7|p-�u �"ߣ�3ۺ]�,��t&cH����iن�MfF{-�×OX�pܥ.�
�v�vl�{�b
ׁ5��1��J�`���ε���k(�7�e��!Ke�M@y�i��;޹�_�`�2�7R�
�����׊C��Ӷ#��ݨ9x_�onpU_>�g��4�.\��B��AѠ�+v�c��W>7չ�i0(�OdO��G�u'�U�q1Q?rU��D\��0�|wJ�`��":�q�����w��Bu��R����"1�b�Vȉ��f:ޱj�dL��1܎�P�����`���B�ǉ>���Kʇ�r�Vӳjrԅ��/�p(��lS���zD+=(*_{��3�������4�ߖ�A�����ڨ�}?2��[L�cPː��}e�O�׹����K��'V��.EwY�ҧY̖t�)��{�@	��NLW���v.��^ �DA��{[=��~yN�03�*�����"BY]�6ޝ]R��Kb@����@S3Z:L)��2P_�o޳[`<L�<W3@�/�>�FL�/�|\:�)

�o�e�.�>iFo���A�Q�b�TG�Ɣ]vA�����9D���yF�ga����nb3cbՕ�ul���KnV�'HW�w�P�>���x�f���Q-0�7	_A@��@3_�&;3��L���UGIlOHj�K�Zh���8]>���`�"�R�8/�k`��;긘���»N(S�]��e(��N�ǊOĲI��^c@	�9���5���)����)����2Eu��I�>�&��~�ߧYɛ.����{Y
�����*K�����P6_�hSV/���S��W�]�8sRVW�2�e��`���ƻy�Ɵ7R�a=,��d��*ͺ��6�x-�f_!����ƇE�&5_�������}�C��!���
��,��Ơ�bC�5g�޿��R�ŵʉ�=������~E��`B��A"�L�bs�Hä᜞�R;67%5H��ns�d��}�f�)!����\�� �!�ͥ������Bz�p�uAR4�c3��Ċ�8�N��m�S�nC�~�QX`g��4�2�ܷ0����^vn�̠����f4�~�����%����LU��o��%2�6b{��cZ*7a��Hk\J�(����=%�5U��,,1�����K����#rzK>�M��v�������!h�p�����Щ��/U >+�5,U;;�B
	~�Jt�*Pͽ�ѱ�~B���J��Znc�� gpHL%�'�r�`ۍlC���%v�~�ݭ ��>�����+�T�y?C�17�}��
Hg�x��6�"���� ��y|�=b*w�N� �bV���T	E�X��J՚U� ��dI�/�� gt~����� ���ֲ�{�����_7 �
�i���xc������fsZ�4:{���l�V��u>�0-(������B��^��Fǖw�.���p�܀v���	^��-d.M/�M_hi�^�@^����m�k�Ƥ�?�+?/i:Ȟx�=���>�.{"�m���2�%��v�m�<�?�x� �!���(7��}��v&����^�K.���XB�&�`�7	tm�@��7��;eT�(���ϖq�9�*]��s�ϱ��2��z�&s���^�a�W�����)��I5m�ܤ�Smlf6�l%������n�w�ێ�Iֲ������PV��	���_�p�ȸ������<�����;?��C�Yd����nd~1�䴝�~�,u�l�,r; �o<�"b�:�����fIޚ����X����qVQ`�B�^�&�f�jK	.'�=2c7w�5}Rn\b��?f3ȸ���*�U��E�ֹL.��F�<Sy�IreN�r�ILC�8��{��\5.���&���Y�7B��"ˋo��)G%���W�.D9jP��NeX(��Ʈ�����H��ި��ؘ�����u�
�tn�M�����ĨА ��T��Z����'�͗4��Ӗ��>.���=T���^�����-�j�e�W������X��R�61s+˒���+�����L��F���� �"��V�u��t�ˣ����a�������F�����nv�ʟ�C'��d��GA��<r�ũ�#2F^�WV���&Sy�g�F)��<r#�}�9��@�I��=ep'�l�|E���[.i0�:����T�P ��K�Lu"wkL�>��]cF�s2��p�����yk�PVu���Bi��<�{j
z�T���D� ��v�^~<k9����TсU���^��8>�t�a��*�3�l��R�!9%�yaf҇]q�����bɏ|4�Q�UJ�wP�0L$�ܗ%���Ay?�c��hJ�l�q�yz��tx]�-3��/=��O�4�n.�³/}䨛��Û2	$��B wi�U�uD�65�,X�E��t6��{U���9�0���G]*�w(`z�c�l��^�R'S��M�A=C�Z ��1�iJ�Ҕ|�dc��rKFv��:�k��o.����MA�����7TJ�P���f�c6x<��11O���3�#sX^m�顔o3�9�ܬ$���l�Df�e�-���R�1��S�K֖�����|�3��g��S�O�7����y�gr�=�'��V��L��>���%�����t0������P�\����};����<����-V-��"�ףEa�O��C]Rc���t����"�W�?|�[��R��?�$&ݼ��8��I�#mGxd�`�	'ۛ�����v�{*N�QR��x���Ќo�2�u�$�	ŽW�(4��N�"N�I����}
!��C�H�h���	�vǬ�9�ƴۋ^FXu�.��gT����Z�ETdf�KU�~{�R�j�
��"�{'�]z��G��a ��*�5;�Ya����7D;#����
�0#�D��)@�uVMײ�GlB;;���d.G�WUu�=�d��l����a��8���O��=�@���\�Hl��}��k���� e��(����R��vT�[n�Q_|�@����5h��}�=3�y����� _��(	���Sy��Uo��S�/e����`�6]��G�v�M��+3~;rzxp���Φ|��%�D��1A��5^%�f "��i��(0>���P���ڛ��]�җ�JD� i��R��/&���L�cm6�\�a<�ruڹ��j`���k?�)P�0-f�����*P�8rP���"�5(�C�
�����G��N� >�t$5x�u-���p���7��}RXG�TB����f�������E��-�����<���J~�T�.h�0x��l���$�Ẁ jbh�&�"�|�W��� [N�/��@��Ä́�_�
�����_���[E(���?�t�s7i����n�X�l~��˙�>����s=_\݋�ՕtPy;�وO3c���L�Q)�\�]*���J֛ӓ8a��F�����{?��E��p%�w9r���9�BS�2�z�ꧼ�Z�.ˣN���Tܮ��QNO��7ű�����t4�(��q������8\i`�b��� S!�OH3���F����4���Qb�189�3�3���b9�tY�����ڪ~
X6񌪂�)�n\��bwO�W���S\�����������@�R����!���T�S5�?$Ҳ��ʙ�c�(<�=b���sK�)�T�sa�J(�ڷ����ҚL������x6�,!����U�ME�'6������X��\uISxR��p�uیvf��JYj-��2�.�?v�	�:�3��1��w#۔٪�`*~��d��H��&��i����M5�	�eE;F2���y&�ƻ�����xt�K�ރcS39&m��Э�D����f�>����6�Z��lǿw�|х�;)���z&U��G�މ�Y�*�z2��|&���������`���/��&Ӳ�+��7;���_Hؒ�/�9�^�S��XB?yW9 i-����ۨq7[邥�=�p�m��*�׏ȡG����ͬ�O;}%&���fB�&�c�&�g��#�����Ɋ�����ɇ(w���P�� X�E����Ã�9CW���?��enݐ���~�4�-\�Q_��fAa��E�g꣤o,H��y�����F ۜ1M1̼�i;���I�$��B�p
��C9�R�?gV���	^b��H������V�����v�r��&����%��NW���4���,�v|�Kr��xg/���A�5[�"�CRg[��͈�co��=���Ϗ	�m��{G��F������gC�n��]/�h��=W��B\�9I�/��η�xZD��&�'{�PL��>-�����K=�Xq�	t����΁�ĳ����T�^�:�0ޔh���S���/��.m ��,��3$�$_�N`h�sz��ZY��Sf�Qa���(���!̛�9��6,��N����P�L��;�JƁv9����╋F�?Dc���^�f�mGꊦ*�n�"�ܡ?�q��Zz�����S�/�o�c�_l=��t��E]$QfV;?��,34q���>	��ï�`�Q���z�$nd��v`pZPpE���ʋW���%��������j�����[���?n��n�HA����h�'��,.X���n��g� �][�p���V�a��K����G/��lXq)u1h/k��O�AEb��̷y�\[�ǮO��4V\Z�g�i���T�������?���zm��n�f��u��8͹� ��П��@����K��PV�cy?�S?���[WR)�	2��@KJC��A�\#?f��
�/O��Fj��3����?�(���I'mYKh�2e�������L�{|Z���`�g�-�|��T�~���n4 5Ѽur�$q9��h@�����4��u��q���t���C��㹒���5��*�#G�������V|W��ϏPfL�����Ze��C��o�Y-w�Z�#
Ր�����'3���xO�y��҅��FK��X�х�ư�PV�c�f�p�6�V���v�3��?cG8�8%�P~A�Y�����$���*��-��c�Cn�'W}AH�b�6o-���P����������&߆���"=�O�r�	�πF멗�JA��^8wϷ�w@'湕EV��r��+���`�sk*=�ҀG*����u�	�1 ?ãx�f*�e۩��wM������"��t�&M��$����KB����zWG	�m^�I�K�+�`��Ra�����,�[��@r�E����o��ݽ�20�����&X^b��M3�*�H���0��M ݀�ѩQ3���=���:���5ޝ�cEqJ�&�C�����)��X$�F�N|��y�?�ME�rP�y_k�V텆�.��%�2/]Nv�$kZ�Gn���Y�5��h˞���l�R���E֚?���.��UC�_�f&QV���"n�w�x� @Q��5`A�%=�܀���4y�=�(`~ҷ�7_���v��S{�s2(V�ii'��96�U9`���Z����;w+ɺ�c�C���D���p2V��$mJ�	4�؏c�+���^~k�����tU7hx��p����n��ു�ۿx�I���՝f/��>;+P)�m�`�ϕ$�8X����rN��"X8���4iS�xP��������4k2��iB��7S��������.(�eU��j�7�.y��3:]dx�K�%įӹ�o[�D�e�5YW8v\�����������;I�n�s)?����rj��Z��	lW�-���N���/�x��	��B�&����u2s���ђO|e��<�^�?�C�}�	m�Y���
`���,���"���5EBBk�6`YL���2?gcЪ1�Go��X�ѧo�gb�[��
�i�hxt�̈́4-'�1���b�zl��R9/s�C���Ğ����<�0�N�WV-5I������[�
�I���2?�6V��n�qn�~���P~J^���@����CvTԁ�q"�c��;d�]މT�|X1������1�}�B�Yӱ�|=x�8P�|�<\����{.'���S,TwãN?Ũ-;�x-��5)�����7�44>;�uW`@1۾+�@�?�^�gsf�K��8��\���*�m��-m�������6=�	��_L�/�X��F�=l�h��Nݢ��k��ԛ��H�^�p���s��xcުu�k	��IC�萩�Ɉ[#95uK-ӹ7��6ގ	�E=�_Eal_<j�8v;)'�]_J�oH�̡����S�Y/7,q��vtp�֐07��'4X�?/t��ΰ����0����I��8������G>0�k�[��/O�,�TɊ	ғO*6�b>�$H'A6Yê�Z�YX5RE2#��A�zV�v��%���Լ|@i��=���8kn�'�Q�tZ`L�=��3�'���k�M�Td�R����g����:�>ْݕe�Q�4�y����R��1Z*������"x�雠O�ϱȻY^"j�5�K/ړ[�۰
Z�m����/<
 ���iV�=""�6� �ъ�`���?��SLuy�g��h�<Ք6��487�4�9|~c�N���
�%�����Z��&��u�nh>`2��*�9��hUAD(���c�?��c�4�S���=ƛw��LJ�|Av'�[2�Q���<�Ū�}��� RB#��bN�ua������ۜ���G�GL�{&2X�n��~<�'VE!�Z����g��G+�k,�|��Ι=�&'s%��+��V�ir�Uݲ�����ߖ���7�ϔ�=Jw�9lU��]���U��H�������f?oܼB�S��e�4�dۗ��L�-wj�Y���bo�F��Q�4�M_&�Z�x�M�Y�#x/��ՠ��!�es8�(�w�9�r7�LN瑳�2�37�4�J6�XS�$<�-�th�t��t��2���E[Ѭ�Y�D ��;XŐˏ���n�v�J�`$���e�x�[���Z
�Q���ň���Ȣ��;�:$Pn^�$ '�43���hb��yF���µbczE�p|.$�?�G�uT{K�� �^�,?P���Qo�$���*yD�*��ކzt>"�H��3�-��./��\N=V</���l�s�&��.1wv�� ����b��3{L�>�r�ۑ�������,/��P�z�w�7�m�$G��,�Z�/QI.��������-*ڷe�f�r��5�<��c>�[�2�z���;/$��-���J�=iN4��-N��%K��\��OC���R�U������𖛹�a�El�-���.Vlė�&��y��'�+�؋������Q�#����BN�w���X����uT���_j;�4-
�k�5�����o���e�U ��MB��I�\�H<��ȳ��Wïou�̌4�{Z0'�U��@�#�UX�}�e���\���"���6�O���%S��F2�gs�9�/��}�/h���e��,��u�QӜ}ο�/PK   ���Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   ��Xք|� t� /   images/83f16691-8d82-4f83-89df-fbd07d8206a1.png$YuT[��R��ww-w�`�%xp�b-���P��.��݊��-���#'9{���;3��<�j*�h�D�   M^N
 �:  0`D����0��/x+qeq �.��� �,o#)��
����������c�b� �"r4<AI�"��+�uiv� T�U������� �`Ll���pdm\<�l9����r9�{��V��zQZ��o�5��\]^�,�tg�N{�`ba�%��!B�+�q�r�c]��xr;��G�V� �k8o/�Z�W�G ,�i��{d�-�]�N@� ء�>F��F�4Gq���Z�sd@2 `��+A����-/��R��A X)$�@�� 2di`�: &Z߀,�����*1*6��j�@�f.Y��� �XP<��	 0C�e@� I�3G���1׳Sa��*�H�JS���mM�I�y{��G��oW'aJ��i�t@���E�#w�4�
 =����,|t�{dylw�{���ڑJ��f�_g4,< Se�j���p	�i�ֽR�X�Xo?r�#��!��y����*F�[�6*DJ���rIkV�ű%�ƽ������u�k�s�X��(诳��G50�x^������HH��X��=�:��PD���w0A�r,e�4��<�/R�'�*T�W��cӄ]��/�(tМ@���5�%�i����  $�<ŉ1� �Ҋ���B��d�aD @*�S��G�>ܪ^��>��^XS)1T�^!L	��@��T�O���+�M�pD�X����}��юw���; ���v�"���"�R
�c�ŮPM#d��S���$S���S���VH�&�Q߲��
��=ǯ�RpE�Fv�r&�W�[�uk+''��w�u��0L-��5�	6��*����"c�����ѫ��a�& "�|�!�W;�L
���#��5�B���
Ĺ@4
���/RI��^P7b�#� s��S%��6��`?z�	�Ńd��~Q�Q��ѣ�'�Ѡ�%� S��sɣ�C���X�5�E�0m������Ƕ��(�Z�1�U_�Zp�����
i����
����%y\�?ԧ*r������{��k�U��g�Ne�KN�-�̴��y�f?ukG�"�N��69�xz|��--hDΌ����Oe�-��3�J?̧e�jr,sgX�c�;j���0��%�c��h������r�]����Y��Qi��W*�ՠ�_���_�XA��Q�W=�Ʃͨu���F����+�����沸I,�hÝ�@ҕ���.�<>�{�UҐt�aYe�`�s�<�>\�s-���0M9�6���U��n�j	�����u��]�\�_��]�;�����>�#�󵫷����Ϝ�̃ϽO�����O7ge����]-]͒�s� ���������@�mZg��w˱&����f��[�~�Y��z�XV9��U�lYl@�L�l�֋�����!����n���,U+Uc��ِ\�����ט���!�(���ԵT߉�ʩU��"������U�K�,��K:vj�:Y�Y�Y���,�G��6�n�㽆�����E�¥��?���̐N�`�.}q�����>�a��y^��3P1X1p�cElU��s�KP�?���F�a_Y��3�rH��}�i��(�#k�j��9)<�W��̖E<f8 |%�����<��S�U��n�a�k��E�ڐM���a?�>���5��DPD��y�NdX6�'/����j[����?���k�˗牿q�=�޷�7*L`�`a��}k�����g��|����UO	M��%ɱ����	̽aŒ9�7����G��1I�D��:�����X��t:ٌ�#k�Jn�)�������ۙz������RՁ�UW�M\Etۗu�f�*[;��"�5��G�7��G�4l7�ˈ���A�}W�c�L��L�T7p��Fa����D���.�n���t�z�� 
	5vB��2eR���U��B���V�ģ�?�7��I>[��ʸs#���>%�Q�)kK-mUͬ:��
$g'g�lR��9ZZT-�������ǉ�����\����B�f���j��J���^���^�r]rz�ۖ�Ξ�Q���v�ת��6��z���P�Hw�SGix�q�ͽl���&�'�S��큀Z���������I��:<)�cտ���x�)�ZW�i���L)�UNU�Տ�2�G{:*Ƌ����kk[
-��r���U�=5
]��?C�Ѡ�71����
[n>���S�S�Sp�������U�|E|r'��B+[�W�֖z6=�ޡ��}ٺJ��lb�ҁtI��;����GdF��s��*�:������?�W�n�v5==�H�@�29A�ì@ǵ��L�&'=&�~��>��R߯�j'�S�-���r��s�=�U�E���]W'�E9�F���-o�W��`��8���ᛧ��I�e�e�9*���J�Cu�.+ə\Q�_J-�cw[�q�םN����i[���²�Nw�j��-&.u���~+����x��]t]~\f3���� nq��$i�m���sI���Ki��'Ϋ�{����g����u��;�&�&3�W�Ha������v�d'e�e�c�r�ɉш�nͧ�v���pf���߼�]+����(΀^W�Q��fz��+�\�*+jG�G�;���oJ_���~W�W��#]��b���f��#e?UD�}���?߽��~�y�`9�2 �C  ��C�' �; pf � N���B����t] ���>0)��� ��y)qM�싿�٤c�eQ�X	V�@��E`e����W�d`ۀG�'B�����@+���#t�����^n;������K��K������?PE��E�����Y�\Aw۱D��
��yw���؟>��<���<[MFp��ZC�#�L��(��~2����;��J�q�f/?3������pY/��q��ҽ�3	�
`�=fy��-�Խ���s��(��eF������� Q6���֊|A��߈c�4X}d��gY�տ� ��4�\�s���"8��둀ĝ뾌��� ���:o!��󘇚�]?E?t��Nf��kI������{�X����:w�6��gx�00�׏fǛ��~�X>me�wd`�F�_��s�4I�e�@q��!�9]�m!p�����#���,�Qe6�j��aල�>~Љ��T�[&��X�9&�8h�R�T��E�*Cm������A�!h��P�p�������d�����/�Ͱ��q�$6eBK�����Y��<�Z:�pj�a���(�s�NB�~Z�����tܥCU˺�$�3�0��G�pƩsP"�;het����o�ǭ�_ʐ}�_� �@���t��#��\�$��i/��:"vA�=Rhj�s�0<��`K���3����Z���f2df?��=֑�)��L<X�#߭g��~��PG���
N�>�Z��}q0(��V�qؼ�\��/���>��`~G_�h�����<�+�L���O��+|����,#�v�M�B.�`�Ew�X��Y�2������*t�>� 󦒊���#W�y���/��{�/A{"��-6���etr����LfH,�q�������V
vD���:0{�3��4�ei��H �g�w�O�0��oN��^5�::)�X<�e3��b���A;�Oc^�k��ݟ����DP���G�#1'VF�&aP2v�������'��F�rDA��.Ո]����=�"�cΗSQ�m<�fuܻ.�ʮ�{F����{���Z��(�j�2�#��❻V޴��4�At�Nٽh���'<����{���ނ�`�����5�+q�5�̐
r���5�YR��{	�e��Ҽ_k�z�k��B��U���U��@^٘�Jfd�ERf$cE�_� e<��?���q���(x�l��n�Z��ێ���݊
G���ŔP��ԫe��|���eTE1��^�q����)�ĳ��*��p�����^2��_~d��ܰ5��K��j�1�?�1�f���|I��l>.Ui�V ��Ps��}mh�Z�3���\���F`,4:����/�*�!6^�-N�q2j}'*jGHI�7���8r������m�⟋c�;�@����,���ُWo;pB��M�Ju&����׳�dc�#��}AL��6���p�hLX��0>����~y��=��� �����_)�3��l�˴��K4>�D�6�k��׻q��)J%�O	��@�	�ݒm4B/��.C��������K+�Nb�M�!�D֒�B�Mѿ�d����rS'�M���+c�tv~����X�J2^ZS6�Yv4�m� �����ؒ�s����#y�"~Yv�k�#�+��x�	��/�8�!��Zp�X�r����1�g��ŭ�]#���J��e6�'��s���mߍ!ϩPa�8�Du(�+ڐ�B�?���EU����h͆'yW�6���f�,˞�O�Dgi\UrD��3�Y뼙�/3��Ϯ1���:��A4��JY��3|zl�j�ڻ��؃{��a��8�*����<��������@A�7Wn�69"z��!r?�AΔ�F�P>���V��+ c��X�g���a�������D�p9��#�RyoH	�v��9MX7�� �N[�F~���7����/�'k�dy/����bR����PE�G��,R.=y��0�`CX���R&�y���dge��L�W�t�8?�/��ꀡ�������8-��k�o�L=P&"rw\��O,f���j.�}�~OwE���ʣo7�l]��i��:��w���A��ɮ��J��g��y=ő��(j�4?�]����ys��㓿�S.�}�,gT�JFqUu������ 6���X��ٌ�N	^����`��-���.��Z��w�)xlߌ�5�����DՙA$p��D�׆�>s#ǐA�jNe ��\ć�MkPg���G�i�Jd��ɕ�gF�)Ag\�\nk��N�e��w�	�~�9ǶIA8�	�"3 A��u�y�J=\9d�kc�������kd�-W�4Z����U���������b6A�{����o�p�������1s��Tj˓?�.���$�ݠ�%�.�� ��?�Q�GͰQॕI�	�)�w��n�ǫ%�������u�JI8� �9����q���a�f�G��K|����7��A�ui��G��te�������-5�%w�ʳ0��gP�۠J@����8)�1bI?3ؙ �$��J��=LJx	�bL��4�^K#���΃bb#�t��B����]�?�����Y_��e�﹎r�I���|�}�(��yC
(=.��*��O���:��zn�w�f�n~d7|+�\��Yb:)���!��x���W&���֗�"�׼Y����bu�:��c뿢�elu�[�B��ďPU���J1�Ƀ3����D���1]HGl�I1|6������H�MH�jC��p�?�r�.��a�d��f,G^�n}��m�r{����Aך���:���D�Vrzx��b�'���
Դ@c�X {�$Ž\�/�$�(�Бi�k7�Z(���GjG:\"�S�Nҡ�6�W5���;Y�hK+\���
9�π�"��`3%=X�7�*���EX����ӫ�f�c�˰��7׃�W�����	-oi/�ڢ�%��k����������F�O���+�0���"��?u�xr�����P���R7����Vur '�SF`0yJ�? �F$���6��/g�/eG����Щ<� <�Ӳ�5G�U����-���kq��z�r�@͗��g�s3�ʉ#�63j�/­�v&��@=��i�l^�7����;�]5"ϣa�M���*:�`g�&`�Î7���C��kjJ�t>��<c�H�JLT�x���3�e=�ȨdGDZ��1M�|�������y��e�w^���0���}-�TN$�(�P�v]��Ѐ�Au#�ŁU�B�ZC�A�r��UY��MZ�F+å-�_wnE��&�m(G����Ju�_'U��z�y|�kzJ�rU��lҿ_�������*�K�ډ�Q�T���B��-������Օ�	���y/�n��ٷ�W�Q�L	=o��s9H�?�~𧶓êԮ	�j�G���c���]�q_��!o�&Gmz���fP�}B�Kh�S]JǓ`S��E��\�&��Ǧ����72�F�^��s�r�~���X��7���p/��p��嶋�*��xi�w�y��2��!�3�K�g׳�8�ג�8)�f�V�UN��d"���Yu����N��!��#�T:%����)n9������?�㐅`�B1��X����[�B�i�Jw������SYO�]W~s��%��1���.��/�N9��g:�A��1LV��ʖ���;�v������������ě�#���E�S>�9k���!�0����UaAA�8�:�V3_V8,FMO-���U��]�VZ��4�;cJ�.�����icڡ�/�X���5��h$ˊ3W���lΡ�������j��Z�b�%��Ӗg ����P{{G�m�gt��٩�G��:��j��Z	V����0q�}Bfxmy���A����ȸ
� �L�gM�M�BudR�S'����Pr��7%*ƺ�HU��M��4�C ��c�'�~�iǲ9�����葙ղd��oDp+Ls�ɰ�x�����߇( ��;F|�h�/�HDZ���ŐiאC�q}�;C-E�\'���%��))S���B����jY�Y/k3l����J��Y�;G���-��.�/,�7�E��Ɍ�8Zbh�;�"x����p2��"���B��?K������fwM���x�Ō�j�NL�N/N
`c1��N^�X
�`�S��k3�C�aw#h&��䢿3a.�IQ��}�	K:�߇�� �lc��ɐe����%w�{Z�,ę�Û4)�$c���p+�q���%M�/ �;I���Ӂ��b�B��ʘҩ��p�,��Z*3E�ś��qPHfŞ"FR��4���~��Tbgm�Vr��گ���HD�{���Da���VV�	�^^�LMDK��b�>����pa�O��c����S�lBp�7e��u�o<���"Kb�4_c���
�%�LX2�Cf�ͩuu�
%sB�*�cAs[[5ph�zn�C��iVtv������KÆ�~���cf���kg}�6�2�w�N�Us-�{ٮ���n�ܲ�ey1-<Y��;�X*Ӧ �I�r��ÌJ
t�y�q������(�T��p#�Du��ۿ�y�Z��/eA�CשG44�L;�S�ڷ@�/����c��y,��^�#}t��i�Պ��1�L�|qI�z��ql��ra�6�2�do���ǋS��H���K��Z�����*=��Y�cv���
Dd���@��e^)�`�	�d�fabN�I<�Mw���l�%�V�P��P4p�#
��TH"0����X���]�˳��3T���~��j�7j��F��1��<�a~?Q���[7i�ʤ�ʹ���-Q.D����owdmh8�9���*q'Wt2��/�[�&lд�`~h(Q_����&�M6���uJ�A���,�K�M�ʵ��q�vbx
ߛ��04����<y�����nZ��c%�42n�'��1�1�z}K�FKZ��c�Hɛ������ɩ�$ɢɈ���,�)K��2x�
B��7�7�)�`'�	�a����bk��G� -ƺze��R初<K�%���AŦ���x.I����:���<�"��+�yZ���rq���k'�i��8']��s�M�o�2����!�U���8��R)D�����њ#j�o���lf�p��&b�����t�q��o���_Olȥ��U��4��RF�w0ׁ\�wc�����*勤! lI�ȿ,����:Z'�B��a�#~�vr
h9���(���V��["V.(��L�����O���l��|�����:�a�Qؾ��z�n�7w���)��H�1�����m�C����V8kM"/q�9ME���w
y�$��sERZ�Q���lm��:z�J�F]?|Y��I�rx:�F���u�"�/o��)�mv<�2昨"�
�b�����G}1�{�,��]��!�A�+���h��;A�s�d�p鏰�u	襑j���[2tId*|�纘��Q����~)�w���sk	m�J��x=�M{�3*����	X!�Z���VOR�ܞ�W4P�aaާT���?]�w9�_�P,�+!mA�t��cF)ՙm�A��5������mp�C[yhn?��PP���ܙ��`��d���;	Kq3�O�,wf!�$��8���������jg ��b����]p�v���OJ���P͈&˿����iotF2��Eo�Z	@ֺ8/����Y�~���gZ�v͌�'��q�-u��1R �ib����t�`�&�8xgPv�t�p�&����.�|�{=��mIE��$�*p��h+�$��vR�kC�������;�աt�V��k;�J�q���2�����)�Ū���6⠚�W��b�Fe����� ��h�e�IM)&"mm�s��Q�߅�db�~�N�(�,��u#�$~��	���/�Mʆ�3��b�ޡQ�*�48}�H�z8#XtM�� ��RO�6�g������ď�E��UɈp�]�Xp�Uj��/�,����IscU_%�k啎Y. �g���#�(���y�z�G)ef�F��}��S�o�v��|\Y%d_tI�>�c��_��]��~ݴ����(8��f=��ŀ�n������Mr�|�����	@��8�&U����#��ם��l������E[Wʑ{O0tˋ�~ɜ��?�D�������U��&�Y��*��:''KWPEJ��ڙ�]�����E��ʢ+~����)�as&���It�$e�4��!^Ě��&���}��/c�� ^�{#	�jPyQ��<G��ε=��C"�h��q@�Z�c��N�����,�Љ\����
��I��U��w��Z�g���y���z7�<x��F�d9��X�^���-��Rl��=~�K���(������������4u���7����,)�`��S�R�Xd���]���_Dy>����)a"��xv�c�F�Ս$�Z��T�W�'�)��H�_lPF��uR�6p�<ݺs�aFxjI���}�I`���7ᥰ�-b*L��4�{��ɑ$�]� �ұ������kFF=�)�v9$w��J
�𐠵��P��ǶH7s��'{G�p�_���Y�V'cJ � )�\�hp�ZŋxiN�F�S8��1�
��6�Ill����=f!	v�&�V���ou+,w����~¬31��y�u7�4<��31��(�rɸ���UuR�9�lj�JV)��_�M�'��t[��Q�c�K �S��i���\G���C�k���E�"���]+@�2�g��y�-݂Y�M�ʹ��s����˥ǆ���>zޕ�c]o1�[�~^)�կ����,�K%X�f��\mR�D�i��w��v6�-�9�V!��.�'��Y�V��/;�|YY/C��ݴ����T�D�_�u"x�YU�~� A���=����G����?v��h��i(gd��J�B�;~�0\9�P��4x��FA��������8&��+�5WeF]��H�f����{g$��\J���`S���e%MOd�0[��� :|�_,�wS�̒7�$�d��9��l�3��I�k]̣R��m�2��* =��%IX�3��],��}�=�;|S��*��AJ7�!�dK+6��K�,��f�|r�'z�]i�8��:5���(r�u�tՕ<S(��U�v�7G�m�S�0�x�g`۱-�������͟�U��|�S=���z�i�?K��������t
�.�)�x��(�oަNW;x�)�[?�LG���_'��ƳP�̧*�;[I���N�}��g��s4���er+�N�X�j�e�Su�����Ք( }�P*�v���Iݡ��V
�ģ�$R\�|��Lu��f|�T_�|6�w��:n�K.8��Z����ƞ�%�i�L�N�ܹ���h͔%ڊ�de�s��{�������~L�D�ժÏa[+"�*�^�_�g};3�7�!��������A�N,t&{�1U`G��1�0�1�TF"�>>X�[����C$�%	R�P�=~r�i��V��Q��P˄&�{ۨ�~����f����eM�YWyi8<4T.����{���S;�cm|]R5'J6}�t���YǢ�0��Ⱥ��:2h��DY[����gb�'�(������y�$b�{i�5��u��[cǮP��[ƶu�s�؍Rh��_����)��m]�1��qUl��_g�B������?h��&S֫���$i��a����f~*?$�"�<arb��^�?3�X���`͚�+�a���E��&wt0��J��V�/U��ڸRϧ���E��'G�"�:c��1����������
��fb�Q\�C��ד�������挨J^cϨu�9�o�{�c%@y)|���G�J�ޡ�6ʍ��2���j���<1��ò����������q��CX*�RYC��������zQ��lm=!8�o����,n���g.}���C���e@�n�P���f� P��CG��I>�&��TY�	���@1���8����]"&Ь�4�7[U�$#=�)x<�м��lXg��;�D���a��7xTo��~{߃��~a�1�o����L֢g�]F�`I]�+���dgbD����j 帼�Bb�,�ח��k��n߹t�]dꃳ���9�X�]=~6K�?<2�<ad�͎�IҿD�T����8>@��Z��.�4��2Y�r��6�Xp6�j."���YD�\n�U�?�YՏ��5��.�T*�b�������-�DK�b�+a����^k��`���#y���3}h�k!F�V������$6+#ń�?�i���^�*!��a�,��3�l;5ҏ�^K^-B�E0;��d\��ުr�:�Q�N�g��s�ѷsМM�� 7��4�>L�oL��N���Ug���>ψ��C�3?��:zH'�}3��~�Z�6KN6P�	�Ibw��C�:ޖ����g;i��P[�T��"��,�F<= ��D����,�,΋Y��;fqԶ.��6�=�������~[oW��q�1Y���Iö�N�UxXk��2�n�u�s���j',������zQ�ܲ��S�F�n�I���-%ן����D5W���]�F��ƨ�sK�Y8̭*�|�nv�Ǧ��n���6P����W��%A��Q���݆v�G�7K�K����9Q<� e���|�R��D��=��Յ�ųT��%���I�����	>��r���j�a�f���P�ܰ�H��8��X��\�U&dWga��S�2��)m��Q�*\�()J4�T���g|n�
��u�n@}h�Y�1��ۚ1��m�l�D�[���Ox��&�Ռ����J2�"R �@�̬�[:�ZR�^,LN3�_��d�7K߳H�\҈ ]�
ʘ��5��}��k�S��㍨��9��}yQ�.��E�ȊR:sU������� 	3�N��p�uǽ��Q@���&��BCH3"e���j~�X�9^/M��c�4�Fpb�0��2I����/XD�ǽ}ʝ�8�dt��O���Ö́�.�fX/17�Tԥ��WK5)4��@�y����[š)�yት!e������?ۛ=)ST#j�.Y-+��mM������V���zj��e�1Ln-�i�̾�M�O�cj/=�>�_�%����,�F�����N>1���єl?��O��t[B�{�ڪp�҆Ę*��~�ac1��5�U�?�s:�(�Q*�'	%�e��%�8���(�i{��i_�y���6=2~����e�|���f��o�VΌ�U��<!J���X��v	S��=+�8��Tf��m�ה���MnR%-�-���8Y�+����a��@��F�D��HLX{�%�eJ}l���`/��PZ�X^y_vN��"LޙpM�/�Ɩs��ƒ�<#��I��.��]�ι�}�w}�I�7��ҵOge1=�j@���o}1�����޻x�£H��~y>���2�3�2{m���5�=!������"C���T�V����W�E�W����w�pM����T�ĉ��#C$$u!�tO��u�]����T���♺\x|h.Ѱ�0��}�TY�+���9૩�����Ѩ���c� q���R�S`J���nF���q�!�M>��C�����S���N����;UI�7���.
a�zǴ}���K՝��j�X������R�'�� �,F|�:�<k0��#����O�m�x쐨���;�8�������"ߨ�`��Ds��ER���.*���7$cϫNH�&�-#Ҧ)��U/��,��a�HSJ 
~�(t��@j�V�5���^�m�h�7��D]��uc����p?�2�$�)�d�䗑4�h`-ܬ |)�&� �E0b��&����V��1$0!k���H�=_7$�I���E�_R��9���|�Oy���>mV��T�y��Ȁ����s�!�R�k����H+�T5k�9 f�"VU�\���u��k6�J���Y`��?L��J�\�a)�VА�_=���QoX*�:��/9L���c�U�\��d6A"��e�oq���cb�e9C(z���$����|.��z�dO�/����=`0�CP�=����	 H.׆ 2V,��C��)�$LB�"b�ي&6�'EG��Q2�U�A7p=r1M��:P����q����C�f�p@�����I���\a��ZS8�;�%�nr5&�
m��NFY�Ps�!��N��ˊ��Cn�/��E��hMz1M�e..�Hr�P�Ӡ#��.����+�y�? ��<*�ٛK O�S;�E��������R�G�#��L|��/Bk[�K�I+�������[�V���Ͻ�2�O{~Μ�
�mէLW�	m�<t����u�|��>"�to����5�������6��eF���4��9DU#2"v�u����*�3=���+��.{��O�(�f O	W]#���I�@��껍���8T<��t���.�(͖�ef8�X�˖���O=�<_��Z2`���8�OL/�J���R�4�Ц������(�j��}�W����y�}�-(�X���_W�5���,������\S�*U��>;�ܚv
��p��[5���\��%�^��΀�K��<��J�+�*�*~h��%�Zn8eF��	�ˀ��?��\u�5hw�h�]�<>�㜝w��>\JB$�FEE2Y]���1y\�?[�g�p<L��7~�j�<�$S��<�ۢ�oT�X�ܴ|�ͷ��i�@��p�I�۝}H"��H�ED^�J!��*j���O��`ss�"�C�>�i��?Y��9.2�~�����<{aQk�->�GQv|�����;#Sѐ�����ל����otr����]�x��1A1�ז�B��}�r2k�p�E �=!1��ސ�JjGdaz�4[d�y�zw�f�ahh�`���[b��/H�"��fY�2���ϑSb C�q������m�q	��t{��^�d����{��(������'F�1e���P�1�;:�������� 3���63�L����?�;���##+�`�E�
@~��Q��� �z��Lwt㌡(��.�NT�,�
��t���_�ޭp;���ݽ��� ޙ�Jm���YfɒÕw��E�������0Q�N���X3)���b�n�?�a�&�ۏD��u`���Bu���ԨHM��xQ��]�Y�X*>�"榍�"�[iM�j��˗����on�X�%�\�,�}Y Z��cq���8#�Pu����kǒLfm�Ɲ\���û�E���y'�4��-p�%4Ed��	�5�.�dӤr(���R��6fxC��jl|�e�+\��:�e�m����;u����w����""A���U��O�[Z�WeD_��v�g֚��B���yg��B�L�0qOX<����jCu��i���A#1MJw�.MO�T��42�{�J��kc1�IPP0�($q�tvN���Z�b��q|�Q#��{8�Lؕ�u�T)���55q���}�:�ں�/>�%=�Ed�����Y,m��T���z�PУ�������D���'���?k��������)M�A�M�8�u���r����\ q5��?�w��j��=�?��:�l2���!��g���&E�@��sw��*����s�����eu�x�nʧ=�Wv��R^�W�Jq�g/�D����l��*O)����Ù%Q����E9������tQ�2��sx�l}��!�H������'!�=�7��K�(����Y4��>3�1+���ߧ�׌�B�Ǆ�����kRS�)�:z�lD[m?VoW��H�v7m�v>��#��x����a_$�ç%��%P#�����/���>s��#�����&�����t�.1ܑw��Z<*P�8P�.��ޞ�}X��Z��X��r�/�΂n��|�@���B!ǌ��Ӄ���Z�L}}����rm[�L�i|g�#%�yB�A�F��""�&������I�:�V*н�ICa -8c>8KAst�%e�U�[F��B�x'e8%�K������W���n�/�
�I�܅�p�MD�4��M���UU�z����4�h���� YY,໎��\t�$�
~��4 X��	0�pt9��8CGU�p ��nP �Z9�F�p=��i���iT�m�}����,:�RA[ղS"����`�߆;aj�i���'� ��u��&A��Ɣ��DP������{�������_�	�X��{5���#���8��I���{^���������Zͪg���GE�Ylw<ԡ`�Rd��3���&Ʊ��J�R��P���l�,���h��{o�-��q�w���ۉCAqD�2�?�]@$�m�|ѱm+�q��fbP#�X^g���8�z�q׮j�e&f��S�Kׇ2�e��!~�$.$���w��#;����>���I�Tw�[@�R_��b�L�U���ys�)�>��һ̴�g2�c�e��-����y&f�ټ����B����c�k����c�ven�;���Xi�)n"(cP߁�E�&>"�m��P�V�|�`�����k��oA����=������_d�j�'�eFd��1@l{�􃵪��������=J&'��ti'���χ.�{���l��澾�3w�li2�	�ÇT@.K�:�� ��Fq�����{��3H����ːuu
h�Nin7���]I"�}0����H�W]�O�J�
����m�J�=.�2�,�m���5��#Y0f��&�6.�%�	-ÐVCy�f3��wR�UYE-�u^Ǒ���'����@�ӳ_Gv��Ä[O�m���nN�}nqQYM.��f~bp�`N�u���qC�Q�8�\Bz��N/�ge�`	�\��[JZS�=o�c�4�H���$��7}J�E��^`��~Ho��3^D��DGGc��>���	���v��j�;�A���D	[��=_ŗVއ+��,�;\��t�ar������6�"<�'��I�L�^ �)�!������zcL<#M[���p��^_�X��!<UxdŽ��te�b_�on����7�����輪��L�{�����C��&��S<uƍ���&̜��p%n��^w��㊒��+��*k�>{}���r�^ў���}���P?U���s��U�+_5����J�׵���n(_'+I5$.7JHi�]��z/��U{�q��5L�466�\`a�k&��i�w���˹TmZ����ꩣn}D�&z1�0�xg��4����Ύd&i��f�N��L��	6���հ{r�p�,!���y�ғBX^8�7�E�� �'2R��q<:�O���KX�(�)b͘�Ϊ�l��̇_`�G�O§ld�g�"V����6'}����]����j��8������2�ڢ#�f��^޻K����_�4�N��Ÿ�(�nxf��`"J���wl�p��üzl���e��>�jP˻G� �m�ہ$�-!2����i�<Pr�@��R���"8�*Y��h�L�c��"ܥp��#��Tw�#]t$�߭�!Z]��@����_q��R{����j�Io�6xO�Y��(�IpL:�G�ҋ�R�ʠ�������Yڑ��e�\��a�$@�[kH���b��s��/>�ueF�&�v�%�������tS���fel�	�����R�p�^f�I��y0T�a��y�6���;b$�>�GJ�1Kj��2���z�����4�5c��'C�������i�����kpw_\����Np��=ww���.��%�w��sf����z��T�+#1rfeT���v<(%'��ۘ��G���G�,%[�z%\�F�3��PTԡE��#�@F�dRJ5��9�6�w��YT���\O���Qܾ���ثL:ya�㽴`ɂ�^���VO���2���L����h�sG�K�UA)��1��n��"��2i�c����׀:?б�e)��L���*F����Gx�qZV����������n�_����_ս���8�(�dGcg�Q�B�6&�,ɳS��cW��:����)?Ԯ�bѕ����h�f�:����N��c���،��p�Sfe�.א�|�"jIB�i`q�$�Oj��[-�?��=�1�y�֤7���9�Z��#��f^;��Y$�;O#o�w�Ő�*� ����8�Xغ��Q?�O�&tA�e�����Q�k��ő)�&����u|$����EkO;O9I��50U�Q�뚴�z�T��]��W��"0�ܿ!4����׵0�^k�W0����e*EjY]<:���3,j'� �޳��6F���C��v�P!�YÏouG��p\��*4�Rv�8%�*X\�Z)x/

\f/�`�Mغ�J���i���e������]i��I��~�w��k�3��Q�����F⢟�v�ER]+�b��gR���k m�\ ��h����(��?��_f����73�0}�21,���}��1ザ��.A2�M$��n�9C/��/jY��@�&�!�A54pj�5�k�R��fK���D���K"	I/�����'Y�O��rAz!���#�r�~��p�����pR��aV�����S�8$ 
@P��s�0�		�&��zR�lS+��� 7M"����gg�TOF���q��D`��A.�l*����yhO��(�	ȌVmݕ��U%t�U��O�<韔8G��������й$��JqJBG)��%�x�4{��j
,�ʥ����?��xu��6a`B��h1�U��U�)Fb��䋏���`V�R�����q~�����'����:���8��ܼ���DXdbkj?�;�ϊ������(d�O@aT�/4��������j�К�$Ӡ� b��6^Μb��2�y�%�N�̯摠��Q��7��f��u��6�\�_P�q��D���;�d���q��2�-�����t��;pI��I��;�@�F%� �rX�9�Ӧg���_%����C� 7Y��p����v(Ceȥ�y��iI����w5'z�ܥ��{7���n�ߦ[-�b^^�U/ʪ�@���]�?����n���%��'Eϐt�u��He%lҝ;��Kn##t�6�cg9O�?�X��Z�Ӥ""�2N�
!zO�ZALʥ�x7�%;[��o���MZ\d�T��V����,�E&IDǞ�6��0�#�_(�C���}����X�˖mE@'��R�h�H��)�H;$��V�F�A���?����z,��J&a�jQa;S����qL���+�`���i՜�OP�Q.���D��	QbȖ`E�}����p+�\���U$�Bn��,d�F��[^� ���`�U�b5�gI�"�iGB��������(��ɢ�oR&��\9*�o��>� �����H�pM�*�!Mt���9�үÖ����y�UTd��3�7fNL�}0��e��:�7�9�82�1'��˽s��!ן�`kCUzBng�B>Q�����1�E}"�禍DT��^���u�����u��Lh-S��RC*C�3�h0������6K��8Y���}V���L'�2��i�D�8���iJM�3Eӵ�xGʪC8��B��+lZ�b�#�T��P�ا�� dT�-��)]7��J�,��WRuȪ�n8�R�YO*���U��%G54�: D����	��A�|5������|9:��mY�R� 9v�5=XGU�d�y>;��#~�������hŠ���K�S؂���0��kZ��3��_n�Cz`��i�N�B%����C�va�?д�hS'2��gH�%��4���mj�`��3nٖ�ɭ�ZXtJ[b�.��%-�mfc���*�$�S�UtK&�tǽ�7$�d���o�>��~o�6�������Gf���Q�j�U<�k��ц/���-XH�40�G��Ab�Vp�6m�#Ϻ9�At� �-$z������Oe�n�y^b8yO��w��H�+�'�P�S�3#Vs���l�sBQEI��K�8�=��w5���"�l�@^-$'zYN��5� $9:�ⅰ9i����q��mKM�6�\�e�uh��3�����&���FT��[���h��S����q�q�5�*\���Ĺ ��FF�e���F%��""��"�s�А�Ke3y�U⼵��A~��*x�VY��8d5����Ŗ�r�?���N���w�Y^s}�����b�9Up�o�@ �QK�Y�f��p�b�H�PݹW<�;B��O�*	a�4�?w�L1j8�U��W�`em�p ��Jq��!���\�9�\(I�_a�Sd��m�]�8�,6��<	?E*��n�VFu`+񅃋���4�<����_h����˚�~h�`�Fk��Q(�,b��bM����A�x��X��:;q�1MҐ˳p���������*����'B &޸ќk]xܬ�|��%�$;6 ,�VHRf2�"��g=�w�m��lR��z^ҫ��+�\�f�'��l>��!r�p.��I�S���K�	����؇����V�],,�q���>��J�C�^��ќ�����Il�32���}�t�sfP\-���K�1\��Ďg��33�adx�ź�L^��[4� ���a����S%9I�d%F����o%�y�H**{�h� E��u����(1�>q`�B�Bћ9�&�h8���R��V�����W�%*� �E�f��T��1>�ߔAVQc��&�ʜX��}.�?����xzE�u	��<?O"���e�[�]8��!;I܃����L�'��21�Q�8ͽr��?gPN���'�r���9z��꛴�ͫT#5kS�`���zs�1�{����ť	��Ck �RŔ���D��J?ҭ�m��11&����}���!��(��7f��}ݍzȟ�O�aQ�4�sb|������F N_;��r�H��P�?���H�,�m)?�\R���=�[l�ԋ��.�?�E\�8����JޡS��tV�o�
�hz�A��ԃ�D�s���f�<,�J$�/=$���@�d0�M�dJ^�C(C��ƀ �M�����؅G�Z�ň!���,�[��6��G��`�mgm��_7���^@A��>{�g���uQc"����G�ܺ��?�]��v�>A�&�ڴ·Q�3��R�8w9�kӆ=G>P�.�K�����E���I�&o�G�m�q��9���Jb[�"��?E���k�c���$��Ƀ�J������̺�-E*KQJ}���BZ�5�FW?�sZ�Xy�>�³Vvź���6n���L<����g��0]Sg���&H3�j�}�L�`&m�J**��$���QՎ`�Z��V����ѯ��H{��D9Ud��Ec�P�P�qZ��򐢐�4���BYƶ������I)ᠡW��A0~�����tޠo%g��4��%��Rʌ��'��2�����b\%�K�֞�a�С�0ols��v,rG����)epU���)���0�Œ-X�I�m=��dīj�����'��$s�QW&�64�`R�I�K��"�|,�6�Œ���F��N��e�B�K�,��f�g�K�&a�3g`�
�d�"��K?)�DS��C)�ZA�gW&TCY�kB�68�0�� �o,<Y#���k�"�4ѭD`��Y�Y�w0t����.t|�K�ICG�b��j�ب�ٺ�����n��G�K��(0�収5{�T��'�#�%��$���(�������W
]a��M���Q��EtH&� 3� ���m���M����m-������2uW;F�����A"H+�.1�c>��ǐ����u��Z����E��ٖ��!�������J�ݍhS�,���Y�P��Jf����G�5��Y0gc����-��G"�߿~���v��Ә�a5��X�5t'�?�S�����uN���'�J�"�#z����(	t��Gjm=�6�����k�K._�.k���4�U�뮌�������^ ��L�pI"�+&����j����.��� {<5�|��m ���ҹ"�5�u'����z{Kg���髂M6:y�����O����i��}����r��8mZB�����AH����<��r�������D�X.��8?���޺+�)>i��䝺�lK��p�JЅ]�Ao�̀ :�O%��RD��k/����Wk��>fd�"#ȅv����`��f���S=�RO�:���l>��S���=	��n�`�zVI�Fr��i+��J�#˺G)�X@dN}&��wއ��M��` Gϰr��12��iBwڍurh9�����i&���k�]xY����u�Xx����	��"�e�}�mZբ�ƥ�s����E.˸3NW���'���,�	C"�������k\��3)��v�P��2[���긄��ҵ��RI������G�j�%������z��czҵ��������Ѣ��'�=1�7�
�>q ��s�������̓#3�e(R���ڇ���������;�\]ȅ�9��3���>\i�g#�m~'�g+�������Y�h~۸�ٽĘο��k���rF�T>�Y,�\�ԕ/�MM�9ƼR��S
��9��~�\�+�D�#�f�׾���k�Iq����NЍ�D�$�� 9���s�Wp�J��76� W$"�Lu�=j
HT�P��|}��x������>�� j�;��PvvN�#M�g�d�8��l\PƵ�XH����	?�GV��?st����yA�ɒ�yF6!d���rS=�5b�a\�yG���� i��b�y���>Z����cTQ�G�����g"�;����v=�י��vV��\;p��f9���Q.)`�3�����q��җi/��7�$Gc2�z�ķ�JT�X�h����C�o������~<>0g� �z�� "���O)	c!�������~���|Y����P\�?��j	��#\qE�D>���5�$��3(��*�sZ�~�W������(\&U�Y�%3~�^-��1**������?oxU�e4�0\m�]<݌ۖ�ؖh�>S�D�Zq��*���hh �bDH�(���^����x��oi���mq�Q�5[C�"C0Ǒ��)��͐|�&������F�	������A�Q��j�8��w^��ǻ������ˉsČ�7�z/U=����N%�T{�h	�p ��'o|q���VIE����{�-c���-ь��z�Ώ{s�����Ek���V0��f�Ӝ`P�.QքJR����(}�D�w����m�J��Q�)��6� &K=VU#FW@���Q���e�����Z;��YT��Ҳ5M�� �|�zx��m��]2R�V�tn�}>N���Dfr.��Kbg��@��T×/�/5����ÒGdK�u�����B����f����J���qe}��;�j�lp;��uf}
�5R�u�Ik�ǰV���c8�M��\�1�������ք�0��5Yݘ�]�$��,�Mgaƀ)��_�N�C;�9D�����F:Ⴊr?����[�+'@�}ůc�[*�\�R-*��;��E%I�.ӷ��!�w "���W|���U�~�����Y��P��6��0����1�2���,1�Լ�Ki1K��0P-�M	�ZcN`!�p$s���b�O?�MO8k,��C�Y5�M9�$�����٫DV���ē�SZ=F?��$�!�
dUb�����\ј[rvI��)F�
��<���~ð��)�.J�n���+y��a��*eR\�]-n��_[����گ��r���4�v��,A���7�簵�d�e�P�M����ĵ�W�/�!�pa���`�(�#���0��15�]�� 7e�Aҽi:�^�`�ڍ��j��jPs�Iˋ4z*��ÙeGZb�-��q$�;��DT��=�Ks"�gUHS�0�|�RXԋ��mV�U�æF("t������W*�ۙ�TMs�>�uuvL[�uI���������Zsf���$���is�2�"z�Y˹���j;�-N�&'�yv�JX�޿�t��U��lR!�9����4$����e֡@D{j�<{�.�G>X�a�%@]���>�u�M-A2�2�i��**%
�f��V,��`��R��}���@"���s�_}��V'�c|����<��M�1{��w��K����@ɇ�.��Y{x]՟��P���}�o�ߗ5a�,�ea���?����?��uI9�^�7��u�� ���C��m��̋�A����4��f���Ě�yinh@��b%!5����Y?Dv0 ��]�8�I�-�tU׶4x�n�'�ul�y��n������nL�Pf� �c�*�j5ޚ�u*�jL=���e�ѣ]NnE�Zg�wK#l��b�ߔ�HT�4�]�5�V�c��aK%�ې�m>/��o�b�{4/M��װ)�#���d�E��h�m���l��K�9^��"K�����k�ш��4��@�5Tmkӗ�1�[�a5����F�g�^�� ��2z����{�mt��ȍ$@
24�U�e��^$�-���I�� ��{�ڰJ �	Ӿ5kj	�z3wD��^*F��g�&F�`E��r���Y�����s��|�syZ���Tۚ4������m~v���h`/�!k������D�±@���	[�4&�x�"/
Ў(v����%<�n��I���Q@G�y�?��T�u�n@����X����}'�:�įEv:�-�S�E~���6Α�!��W�A9`:�70��2S�
�����y�X6T"BE�����kũ��z���r>��@XV��SGk2˰6�֟�؛ױ���[㫇�U����u-�29� ��)+H~h�����ۤ�}T}x���%���~���Yј]�}m�E#�[�H�	ÅS�Q���D�(E$�s�ٍ�"2ޓ�������9W��e�p�-8I���1Y?�����=�s�g9���S���B_�r�����	�8������o����+�:�	�)�w���Y���\��4��y�����
u< �'_k	F%�D��]0�W�HV�"�eB�S��DMlrMaCKw�㗌Lw��T�vd�q9A ��ՂWX��ز<; ����T��qt.*(���W,��	6㘺��>���JxTX��Ux������7��gE�ɝG(+li�����y�4,984 �{E�J�!L��.]��5=��`%�R�>��DO=��}��>u�e�&jJ��P�~.��E(��*|��Z�$�sl.� }b�S#�mxPEp.�.K�kB�Y��Y�7�����C�2rzY`�"\�\I�%i��T��|�}U��娠Ω��U2��1�l_�2k\�U�ߤFKO����A�I]D����X��9�߷y��Z�Ol	�� y��B��J������z@�^�m.���)	���yÙ�W��X�:��B_�]-Dа�d�;�g�����ٙi�%�J�R�˵�;�6�V�;�aA�敋������/�����w7MFe�X���_Hד[�Ӻ��~�,��ʗ�c6����/�sGd���Vz"?
t��XG�tc�&����.�Q��dM[�5��$�r��-���~���O*�I��ܹy�Z��,�Ҥ��p��- %�(���e]�\Ͷ�q�$�Qs$�7���o�+��B]}�Ҵ|3�t���(��?�(�Q;.Z)+���'�twe�)+����Kږp�wN�k�ѵɫ]�q߸�j�'ۃt�nn���頽�3{#�ƽ~e���z[ � L擩P0[ьnju��M$����'�En7ydص��2�l���'fP�⩀�^Mbڍ��G��Ƴ�n�1_8��kz����Wu[tJ�m~��ͦ�@/�u5�w�4T� y��(�1����w�l[B^�K�e�*CZ+����j:�zDM���� 6��6P�����uc����A?���t% �ᗰ�0�~@�)�Hޟ�~��A�3�d��X�>}{#ϙ����ȩ�$�#�jٙx�.#��~R�p �è�V����vD��ȎB,)U��s@_&�5�c�_U�֦a�t�9���4�H�c����=E_�7�&ƨ�!��c?*��V�vLQl�p��=���7[�jL*ad�<c/��0.��Kv��*�Y���ɴ
#�F�/#8:M3�Vr���th���(�*��&��q��߀2����qJ�I�fߊj�C���׶�����g�7i��tzo0$�%�&�(�4����cmv����?�5�yݴ�;B�s*�ty��J��愛M��L�
�	m�9��U��k��������ǐX���>oH�I��d��j��ёcȕ������Ȣ?8�/���>�?�Ǹ��p��Pws����u|y�?�lǧ�~~�����O��Un��_������:��-�#K���+=��j��'��Y@N��� b�%4��kFm�=����E0�0 �2b5/���4�~���^�n��[�즱IW�l}o���2�IE�T�ڎ=H�vo�2
:�j΅j���D4��n����$��u��,�!�N��A�S��P"���� �����ў��:�CfK[���${�0̺!��ZϘ���&��>	��7]P������Af6�5gn�vY��kL�˳�i�Y,w~a�`����Z���������W��A����z��Z.��d�E�u��v ��~Ɖ���T���`�5i����n�f��9WiNB�qd��p��چnf���s��zFG0�1v =��Xt�8fb5�8�`̈́�N�Z����RVpȯ�ۮZ�����91�.�>ٙ��MҜu�>z�<v=yL+�(�O$��4ݟ>�Q,.e�\X�豔�i�$�.g��$�ӗ[ÐpHGQf<�Rf��45� ��i+ӑr?���z���1�M;�˖�����؎�(��)�F�S����L y���d�1�X���y�>E�GՅ�*�l�/�_��[�Hg{ٖ��K���y���l��n_6x9��u�ߖ~-1�0$�F�	�Ley�F�G9� ��6i��v<j��,?M{�n.`*d%p :<E�볈k�g�e^���G��a�h���m��,1���v��0�#w��5�]P�G�� i\y���*t�(����2<B��n-����V'�P�
U��؝����������g6�J��1�v��i�Q��D�I]l�<�0���Z��rg��w�	Z�J)��nɟ��U�;��C>��C� ���[M�р��aF >"\��7cek�iō�#Ȓ5�����Ѩ�=k�6��;n��;����t�1ՇjƌJn/p�3��b�9��X�q�gt��;k9��U�5r'fuՑHW�[y�x��/F�"��kP��`W��n�b�`�N�:�����-*���"�~'TN����Y�E��G+�T%��1�&vS�b�	SR�6yXV��c�L�_E�v&.>OQH�d*��AF2A�T�l'�7�S�0�ɓyvO8 1�rڴ�}�%�1Z1�JLRG�������[`0���?��~M�#H�3��FA�%G�Ȕ����$���9�w���q&9��ۯ�i�d��o�(�X'���Ж�'�H�﬛:S`ڧ�����d���\�><uS�J�L�?7�#\��#:ekd�N�t:����CQNB�r��TlAyi�[��2�1f�b�,籗�)��h6�ʊ�E�E`X�q�uM�T�F�{�)��f����u݀*<�<���ʪv4�w�ۗL�R8�O+���6r�<�h��짗#~k��yO�W�^%w�?�w�y�J��~�%r�q*�J�z��D��+��{���ݦ��惊^�/Ae�#w�K|���Z*�x�Z5 *7�H`�Ȍ��\9z���^*nj���,�"�ˮ�$=�fT��?�2�7= ���������U�x-�Cg�@Ӭ
z��X��[&������N���5����R�^���c���gZ��Dt�����D�C�C���!><>(��)�V�I���ĖIJ��+�V�qZ�%|��IOV�β0�_2ᮒ�Ib�}�<��B=�1NDٷ��'e4|�F_L���b�0h�$I���+P�L7	b��l�eZjXc/6�ˀ3�Bwj�L=���
W�D�k��L詡�T��&k��{�ao#���恿T%Z�u��Zz��U7�Ǡh��ϴ����I^m��fK�ǉ|"�/���t}=�5�&����$�&(����`M�$�0e�3��'Ƨ4@k�Te��*Y¸�������3���≮�
��i�������yΚ` X��uY�:V���be3�9e�`/��y&2|�2W)��G��j��_����Q,,̨Tk���s��˲4c�����m���NV)�n�%�4#n��A�����=A��71����D�-�(�f�1��z
��p�KsD>�8 �M:�э��R��J��Q�^�l��\?���f�s�+�����҉�دx[��)�X�1eSf����G�1�ڥa��.UN2(�ng�(1'dxR�������-fq+�[�^��,�׃8a��]�(�
hl3�`�a�PgZR�7�bL�5 #,����k�U�Za��ڼ��~$�;5%��E.��H߮�k��L<���3����cx�C�6�L�V�=�u<6���F�5��LA@�1�`��[�f*ڢ�Xh�|�W�/f�W�e󐾹�JY�%��!<�L-��]��E��t~Ir&�3�oؿ �b�峳�KU��"=(Έ!�S�`��{���`F��Q�q��$��wB��upDiy��R5?�������	Wf�aC��NK���!SNڜUu����Ą&�K��_"$Pа?�U������(���D�@W�1iE�?����B$V1����������~���� ��%�HKh���x��s��K��3�-��K��JI��l�zZȌQ�@��K��d|
{�퀔`68f�2��`6�c��
�b� 9F'*�
3�v�*����i,��j�l��ĉ���*[�2�T�s���5�&ĵ��}k,>�p�ۥ���D1���h���K�
��!m�<"�[�a�� ��6c)+�f*5Zz�>I�[�7��:툒p����~�*�m��Q��ӟ��7mA��~���&~k.∴u#S����c��*9�����Q�X�p�B�����6��������>��^���[��B��z�O/v:}Y2x�'%_��?��/bv�'IU��p_�r)I 0Jه|f�y��A�4�e�xz�r%KmcGL��	�G�����0���*&�XZ �ړr������2��Ȼ��U�fQX(F���ܖȓ"�ޑ�O �`%�iT�����07���՘T������Q���U�y>/�z���5�j�l&ED's���z��W��-N�����ƀ�,mdlqR���ꏑ:N�䈊"���R=�UPۀ7�3~ϔ8sk�Y0�e�b5��C��!�"�-��ab��7���J.M�o)y=��-���v{���)�?�{l1��ǽb�:U6�2�n�w��dTJ�/���6�z_�n� ��C{�3qTp�Kc����R�"��cP�%gza�o���)�Ͽ��K�"_"<������"�c?��l���`������fU���{�����?L�	�y����DX���<6���%!�ՀH5A�Ѯ��9���|�0z�`�ޛ`�0���t��௄W���Z[rٯ)�%�H�]�BYɚte�p]j�mף*:�!U���/�I�2���t��(ח����~GՐ����,G���T�����G��S�?�{�P1�[��'�?_�Cg���viB�=.�S�?�6�N��OTn�޻O:��*��k�j�U���f]�����Ob'<Q{Q��V��>2Onx���=,t�%��6�GS[5�M�騿/}Ё�;4Sm���0`��Ԋ7U��E�߿��M�!�]�ol�뿱�E�t�"��f?�'������?˶d�*1�z��B�b	xo�_��ԘIʨ2�:���m�@���	OT��G�	�J*ڌ��� �/����z���;cB[(�޾x��doObF�u�w\�������P>1rZ1��?D��ow�:��8![�3����iB3N�c�o��v�P)"�T�����٪Ԍ��Eȑ�+o$��!��}����� ,��n��~~o���^�`g��t_5|�OrI�_�B/bTڞ�#^�/^��|��k�.��7�b��`���N��#%2:ZO{ƭ���s'�.����K��C�m'L�ǃ����� �7�L����чE��ٯ%+���o�`��x�Ya#r��#T"�){�X�&��x~n^���)V�^���Nʥ:�3쎓���x��ń<��2B�:E\��[�׃
���D�~�۰���Q��7|u������-JέR��'~��no��@�}荌�d�I#/��v�C�3����Uo�V�	UrPReDq>�A	�xO%�����	��)���P??
:�$X��챳�����+�����Fi``@�8��H�Z�U���`	:5n��Ѝ�dH����q�0���[��+�ֻ�e���RÚ��'[I��/��	P�73�Ë�ʷ�J������V�Nb�� ��)�ǔ��׍g݁_�RW5bz-3;_W:������^#g?fB�Q�KJ��N�x��zIE��C�������ڕ8�������	|�0a����������-L��]jHtu�Re�M��#���ݔ]X�nҔҿ@q��c�xO
`_��m6�z�����\"��$;�=�+��H;�c]D��^���Dw�H����.X��r^��+����?(QEϽN�LTv�aТ�B���+�;\I6�n���t=���B�֐�<�OE�`ټ�b�u��>Cͬ*Yi�%�,qd�l�����f�[ٖ�F�*�Τ�9[��F���e��3)��SG_�֐�d"����0)���hkQn��|�O���U�#�?kr��P�O�v��j{o�=�T�הz�a}ʱ�e�z���?	^湸V��v7��wB����n�*R���MNo��
,�B]�f����o��	�3[���*O������m�6ȕ��;��3(�9��v{�o��d!��-�I�E^ws��s(�l��k�Z��P���}�h���;Ul����dI�ս<^����;1��d�H�a�f����z�����м���+X_�/��M������~D_���MT�1�w���Q�^���G��z�����*V+Qb�����e)�	���Hk�d�_�K[xy|n����z�����
��*�����|������X��J�/�����d��GGW��=&�C�v�w�^K_u�˜�ۧH��Q�	���v�����˵ݶKc���B��w7o&�޳��x�L��~ZqV���[G����U�w�C���L1����B����	�pk]�Лs@�ߥ�uz�m�����V�(PO��cf�?����ކ�g�:�G��r?��3�%�����v�F.V :X��-�j�e��/&�z�zd��M��=��(d����������%|�&X�]���9����M�����q�\�����@�#hg0�ƠV��no��O�J_�R4�3fq��n\���H9�۾,3G�c���؃�{$*1�g����+���w7qM��G:��^���v��yr۟J�ߊ�}5p;O+�;qV���ڑB��i�@���i2h�)�����׼�0S�9AM�3���vF����`@�V��`��rrN������@�o��"��G�"�gz�G9��)h�U@Myr�S��^�7E��oB�i8�ON�΅BhC������RI�B�.�V�_��Wu�]*][44w�m�?�;p�C�VK��j\��T�X-�}Ut��I�A�ƯÃ�am)�	G���F�9�S�5{��qbm�������f�^+[k'�suW)()����x��~Lq�9�y�s�nU�x|�!�؄b������jV�ڂ�|��ȟ�t(�w6c��z�|�[�9h�r�K����p_Y�B ���~�x��ŀ�z�O �J���/��7�{��
�J�#C^�`�ɥ��.7E�����;�Z�����Ox�V>>Ox�n ���q������K5��+��,�H���N�������]�L�w��]�Xk�v�8��}�.��x]��B�J�-�oK|G����6&�Z�ǌ���n�燁�A��ZE	À��w�D��ra�VT���f%�,�Ý�N��W :>^A&���5�k���J���T�9�8<>�m6�2��J���1��9^����l`�o�m�'`����{�?0�\���=��[/�2��]>\��ߝ
!�Ӫt�Z���<wQ�����/O_����<$G�:�|��+֛����Z���+1E�#��9=�N�C�N�����+-J�����3>�r�=}f|N��7ɀ������[j��w~7?�b��i�,�K���ޢ��nG�f#B�/y܆�ӔzN������fG��ƃ��$1ޏ"��S1��D�Ot�
9�%���5��Ku�\$nW�f����P�������޿�G#$\V[�'�!t�O���%
v/��L����%W�3�'YV�HA���H��F>��R�SW��tP���s������G�M��P�wv#��&8 ���8��_���v9���n�!~;��X��<��=�_~̦&�0����;�ſ^�Q���|�G&�!�z�JH1��y�mi�[r^!�@�����"�)�8`�88���!�:	����o���v}��{A�R��G;���8F<�����K�#L(ᵃ1םo�̩8���6����9۶�p��Tx���a�Ǳ(���	�m�?�gce�kOn�����ь�)��m6�x`�o?I]���<t}��r�����EL9��ic�*�xm��
p���.����j���G����m�Rh�kO��C��~@R���{~��d�����[��*�"��=��~ex}�(A���C���7C��o>�O�ib$%D��a����i�2�nTx��,�vL�AѽL�3�{��#f
6oH�� ���>{���ڍOb�C<�+}�88�0.�kS�����z�F\Eׯ[�֙�@%��(8���w�v\<7�8W�Z[/�	uu%*"�N�1�$��o�!��2K�V֜/N4m�>��<�_�dee�.�7��Z��]W���ڮ��.]!���+~����/��Q;�'z.5	Ŋ7o�7Pj�������W�R.[׍L�������	�z6�y#��]��[4Y\x��/֘�c3�n�?| .�Sγ
AF:{~�R?�����o)�V�_y��޳�K�X��@.�ܹ�w�&��a����)Zz��r\����f�0�x�[jp�^� �4
=g�@)�eW��ܟ*8 �����NNv�|���?��I�7:)w-\(]lwJ��}{�8�|k29kAj{.}w>��ۀR^]�F�?������2])��'�mk�}�'xcH�uu�Z�������;u��#��K����Y+�B�م�������k�����L������`�|��r�ޚ�zޖ��u�2o�*  ��z`�}Ї��,��t6�����8�x.�7IfT-��9[��X訶��vY��߸��x�k�dyꃵ�|�(/�;��l�[�ʟ�Z�jz<N��/����k�HHץ��P��Eo��+�@=G.��[6�������f�-����ᵍ7¨����$����R�>���l��q��,ޡ��c�IG����uk��x�;шv�|�t=�9��@�?B�ڏ�^�Z.�ޯz|Q����y��I]踊"tH�x��ĭ�{X�t��U��ޞ�nO��<���^��I��f���BW���e�-;XoS�Q�B�$B�*Bc��n�Gŏȝ7�z7�V�kE�m��|88M���֯�]���_n=7F�����W���l�l�n vBBW� .����'#����5H7p�e�>�u�uY�t:��%���)�v{L�r�xZ䶙x��;�/�v��;!��|c�1�=�/˕W��r�V[���S[���-�W%=^�Tȫ�˗�����x�J��7N���ޗ.O?�73��A�9�K�>�����|�t�p�u���>k����1��U![p����x��6��kJ)�P��/�^(�ťw'�k��P
(P
w����|���y����ٙ{g����yNo:���׭L�,)�w1d4t��4�v��d+\�v�q�7-`��d���렍��ޘ�=B/���gl��C`�����X��d^7�а���F���I���^A�ѻa����S[+��xB�DOR����6قG�s�)[��R=��a��>B���o�	CJ1XƖE �rg���R���5��xry���ˈ���'��)���i<rB�/��I'b���f��ϨU�ē�7Er[��|�Q��IT"�ڡt��1�=��Z|SjG�:�T3���OȽ/HI��2�X�|����Ơ�8wOh������G74<|(Z�0[6��?a&$&�퍗��B�R��0%����QͿs�TAQ1�/�k�/!Y�����K�ӖB����P����E4�D����v��=ߚ�m9�r�G�O�9�W�o����?MZ��e�^Ҵ��7��~OMN�[;g�$ޤ�����e�z��Y�6����o���fĕz�wl`�p��<Ga�'�n�p����La�{kF�=7�������b�$�/,�h�uQ�bBMYT}ʡ�)RGg;u�U���0�)�gC	����m9�'o���uX�	���|��]��p_�T鑑�JuV[�3��ɽP���V�����b,!)a�^��D��^�Ҕ鲹��D&�_���1�{{#�'��G�.���B�jW]AA!צp�u�_b{4)M~�1�V��C���� �]��&�!I�I��a��� �����ݝ�"M�^/��?�ê���ʡ�ϼI!���;V?�ԳF���E�
)ƨߚ���-��:��d4�f��g{�-)d����A�k�.ʌ����.��cI�	�Y~K��TUU=KtƋ��>�s���_r�eT�&�_��L���d��-��v� .�|7/�i�2$Q��N���s�B��@�ڰc���;����~�1&�N8������ꎾ��'M%���.8�y�q�խ���&KR������� ������O�wr��DX�W|�R�a;��#��}�3�A�����t,�$�ݝ��Ͻy��E^�"�p��ӓgAq}}ڥ��O����߶pu����t�-�|;���3Z}&�-YZ�yz�2�o��(��*f�A�S�7����#�aaｷ)I~G#e�`�A's-���&"p�i�p��ZR�����}<���vcuk�{0�`)~���>SL��
�*��IT��>5m�P4��IC�W�x?!/�m��90�#�x|�q�����ǚ��w�� �&1��md:E����򂝻�!*貊ڳD��K���V��c��=�U�︻�_�u�q\�z��R���2(���uH��0	x�Lm36�X	jy�3�8+��dG�o�ͻr��!a�+��uv�Eg��Mϩ��g���,���V��rE|�|+�ބ�j����C.�DQ*������h�ܧ߭����\�CoJ�C&ɛs��]|�ȴ�ڡW�ܜ�F�Xgq��b�e(y�����R�'I�t��������,��Up_,��c0@,u��)E|H㷯�������nV�}��!�V�{���ω�_S����@M�t��]�����e҇�|K+�H��I�)ɩo	'�
N�����3!�O�T����h��{�ś��a.��N��Ɂw&���N�E�PA|6�^]csm�t���gF�|/��uT�XH����Eaw������z��9�U�^��]�{�3	W>dv0X���[�U�/��1�#��6��6d�p��˽��mT��@-�}��b�I�[���s{�jB�e_X��_:dU(�\`�)o�G���O��.�<3/��ɪ�E|vH������$�dW77�==��S�u���B�)���z���u�����nd3[)��<���ub�����ٯMoLz�u�	Xh�v�d,�?jkOKR�HY�G{7���Ղt��~�t>�(�������補`��8Ѥ��щ���vM[9��@m�^S���o��O�Z����w���i��_��|�^�ԭ�W������"�e����t
A�*C?F�ZtZ�]v����G�x�e�ӋpY|G�n���:M�zs![��p�'������e!�� �i��w�]ٞ\�S��&�;2��M���ʕ������S�������@)ZLG����鴵�v(Ѭ�EtGܞw#d>�;�uߟ>�̓�R�N�/]D�^=p_]2H�Xa}D껻��%�����,l��E�F�O�{�痄�\��;R�3����t���� ;w'��^M��{]��}>Hv��
6��,)���׊�}!)$��m��~�}z��r�d[�����C~L��oϑ|z�0���sb3|�x�����\c?��?`�/Iݟ:��U,C�}N,���5��XB.�C6	��Y�� ]{׉���4oG��q[�	���G�ο�����p��u��z�XfU�r��K0|H���Z��=��~�/����'�ۏ	��.}$/s�����|-��J�~��.�Z�#��h�;1n>��8����^�rC�HYȞm+�;8{�+X�Q���3>	���������~X��X�v!oU��J�'˔�3�ԕ���6���ɮ~b��@���b��|ҙQ��r*���q��с�q#n�,fw����\�}���w�u2Z�;=� �xO� �s�
KU����>��c��a�P���S�YR���{1���T�Z����Y��9ͳ�˺'��1�{Z�`�% x��d�'�e"�t��4��<���n�����fu�fBז[3ɇ�䳩��n+�������8%	�[�8TK�5_:�nr^��Uɺ�5wfu���V���pӸ�I��^a@��8׀���d᤹O��ظA�}�y��j�l�Mtu���\��"`�{U�3�-�K�!cd�ē�J�aG�Gr�헁�H!ߞ����S�8c�.6�YAK���n�;����Mt\�N�w��m�'�m��~X�s[CoY�'B��}gͲ̌�wa�׉���*����ն"�2�.���r+`	�Ó-LW%O�7�7v-���Fp[kAor��y��n�޷����9���ɦ���K��%��Mݜ� ͣ��|��jC\b�`�;hr��b���˫��F��VT\/��rT_o�9ZȦ
��m�eP~pZuǪB����J���vX��� P_��{a!�|�}y�j?0�O�8j����ĦEm�K9�V�rs�ܠΏeY�.�4���b�7H����=�̹�zLOyW��<�����Q ���	���.6j���|�0�Ui(Ue�䲮P��u����]�K�b��}��`��b���I ��4���lI��|+a�U�����ֱ����n�>"M�O�+S�/��&5밢9�7�nN��l�}�yOZ@>���i�G��Ŝ��=��eT�G�������� �E#��K� , F�wi�{��H���f��s;U�q��Xtb��	tC���j���,� c�s_PPm���~h��B�7����n��U��hAl�#�G���Xz������vKP��/���g-����W�"����l����"��c�Z\�,V�K,�XZTMN���9/պ0�;.ͮ��@7����ї��:k� ���4���>'���yS�ߨJ��Y��];-7䤜�r���O�a{JU����B�0�p&�t�6Y�lLFS]�=vc:Y�V~u�R���=0lڿ0�.K)/�*.�G� m[�!�.4������&�`M�P�|�	���=W#4�s��-N��D
'���Ll/1/�	�Vᶖ�8\V�Ym���m\s�Z �g�F��$��������i�Ke��9u��I�6���s7'^�cH��)UA涊)Tb>u�0�B�.U�"J�AΫu��M�6js���s�U��9/o�{��i�6�To;E�We��n?'=���Ec��g5V��{?��LU��5�\,A@S/�O�͉���hP;g���& |�ѐ[�X�n8Q��mw C��v��r����Y�WoA���|���Q��r�N�(�R�0�'Bk�aLq�,���_���	X� ��-���!~�5��X�_�4尉5Og�A0���>;]M^�x�w��G�u�`3�6�K^A��٩2�gn�XZu����[����ꟘXf��Q�gW�tQ��i�Ç�;�T��}������5\NNI]���c\IRJ�,�^^�yI@=�=�#���Gw �J�Xs��I��^�n�9�?!Q�O��9MJ�v�~�Y��ӗ�����`jz�|��S�}��`�u�6AWWWdd$���ZXM3c�&t_�rgaF)]���+��������&�b�D)w�"S�7֟��0r�D�w�+�@����d�|<2��O}�dMJ��oi)�����7L��xZ�xh)��TUs\5y�$7��U5uɅ��\(�_�+*����rc����S�Ď�U��|	2,~�K��M�"[4�%_�7�--�ǐ[9?=C_6��䋁!�\tJ
�>=�,w��O��4�W��O9���qI�d�4�"ӭ�	~�i�-��'�Xut�y���Ǥc��N\��O�`R�D�H�=� Chޠ3�c�ضO�ݔ�Z$�҇:�򾹹��3�x^�����Ԝ��6�v�rN���c���wA�Á�F�KE��.r.�y�ܼ���@�&3�9f���;�sĆ3*<O�eu���P�<��͠�e�k�gVRz�V&�'�U�\v3^��kr

ߧ�ϱ�[�_S��W$&�d����S�7�[[-��v��6�6J�oc�������3Ѵ~WT���zz�t��yh��طse\/ ��a��^-R�t\�L�񓪲t���^�L��/͊*6+&gVV�4 B~���h4�X�Z�i>�p�Q�{ߐC��Y�urծ�[l�Gķ��)Ք%7џ=G��}s�(_C�}�a!��thar���q�ˢ�R�0+Kg{���Q�86#�3��}B/��}[�J�L��F.�k/�)ǋ� m��X\-n��U#�����s��`a�)ï��-<�]\�M�6�o�U��U%�5H����E���v�	4��h�F.8�2;�w�w�_�g%��%�vmg�����rDh��g' �o��h�y�7�"bpj��|��@ c�L�9b �aI#��T��s�4�ss�ee���!�3�R���KZ��M.`� v̌o9|6��m��l({В���IYm-�RfN�`\�ʬ㘍ŊR��������]�۵@|��P�i*���%�#8�`1ɇ_Y�M���u1%���!�N�]�0�� d��K���ϰ�z|f��5k�P�͌����L�hy��c�$(�CB뭭�$�r�ES�]:3��D��x�� �\lc��vqT$�T��-Ƭ<��
�PEquwA�%���������+����f���ns�xB��nZ����]�I�#�v҉`�����i����	� -Ti##r�u�s��2����S���Z�o���F�7�Sc��ȡ!��6�,��૎JM(nM� ����#E!1�  炤�Q�xhPۆ��������YTly�=e�� 0����.K�)�#��ߔ�y���O�l�n'�tu�P��� A`%`iQ��_��7̵F�*�L&���C�[S�}���J�ol����=?����{C�
��OO�����uH�ќ:W0X^�[� �u=��V�ۢ�74�Ɔ��+�/#��J�����ևzUF?��r�S�/�P�F{C��������Jgr�&�bQ���B�Z4͓G�@ù�.���h��+��.��ѿ���II{G��9`-s� *
�����*r�;;�!��?��2���p��k"`�ڲ���|/W)�H8��u���ʽ,2�d�S���c������?�Ye�-�$����̹q5�Zr	��Yh)�-��c�-r�$�om�i_���L��[C�OϞس d]���퍺��H�*3zg�P4������k+��9!Z����f��:�Lߎ�\^��[*��_L�{��`�)ȠۅJ
>#a'!�ŖnE)����4Ĝ�wE�!���j�5L��%�=/��g����V� �y���ޓ9�gl,�[���I�2��p�PH͈5��~	���F@���/�A���㏸����]��׋:��~8�KHF�Ѽ ���r����'���I��8C���ill��Ĩ�GGG�����Gb�|R��қ�xk��ITLRRHmb�O�S߳�/��*���j��0�B&&�K��?s����uUU���:e���y�z՞ӷ�d�a* �$~��@�\Y���n�Nd߮!���i���!:%�:��z[�
���;��7J�{d.m�
_-!n��Ԝ�|u?v?�A��S�L���O��N\�($ޕ�ad��{�Ss���t�Pu/~U��o3�ul����ԄZ�1܋e��.<q@?�s/�>B���뫼���Z�>���T��W�>�,u�M%���g��q���#?O�uBTT7�i���<�$�'+V��hi�D�.�o	�i̜����oO/�h���[�I��L��®��,�^��
..��?�v���l��iq�����C�͂�͡**���R�+��'�6��+Z���WA�𣊦'�y��
��}��~��Q��:�u]i���0�wX�Z��|���r����*�'��m��~Ry�n$P
�|�p ��e:y7���@81�x�#�H�u~��
|n�6�Z����gC�_���f?H��[e�Q�2�,�[�����������b��%��gt|����朆<?�����r��˜�/)�&42;WV��X���.-��5,�^��������g����>�w]����~�֢�4�J�*�h�F����?=	��挦��Ia�B�A��-�/	�?�<u[(rD�4���U����5�3B��٣�
���f�� H4�.�]�hy/�/C�ŞBQP6��[o"�~Nw�]��n~
�_��zWS��.wmVt���%��=��+�GH8l����&.BK �	j����ʗB�$�﷒������!��M�6����$��6�/C����0ġ�Al�.��G��=���b"�
�#��������~=�ݝ��i��~�� ��tG )�B����ٗ���1��ih����;���_$�X�6�8*�F�q�x���wʚ������� �Sٖi����q���M��A�1`��xM=�o����tyX����}UPܦk��d�����e��pP[��Yz��3c���^�j}�T��7�3���#�������!�W�\���<��8��w�^�g��������)"���b�"H�Wz�}O��nec��\y�����dϬQ�(!	�%۵s�+�6�=���Lt~Gl�k�7�D��?	�W:J�-J+�*m&�]�4^ %�ٰ"�>>ke'�E���=�f
,_ z���|-m��.�xWp{�2�M����J��?*I�ؿ�<���@�d��]���_�&��Ͻ�f/k����\o0z�ڗ�q1�.�WjN*4��_�O�O�|��o}�����g��%�?9�7�r�l�T�OeeáN?|�W8�!8��Q����n��CPh�W��ʠ��k�S��n�x� ���������V��df�2�q�L��a�,���������֝p~W&�>-$)�xq��nc]��/�>��T3�nN� �|Q�!��|)�G�b��&	��HM�:����70�*����͵p���7�9��[8��/T�\����C � Y���f�����z�)o�A3�sv����n|(�U���&Ǥ0�B�:�;���j���*J����j�z���.`�Z�7�)2�	�O��"a.�kj�AgS�^�
�e�-���2��
2�|���p���;У�	H�M
f� 
*�ŉ-Yx�2�ʙ�T1�#,j���p~;�x{{g�G�^�Х�a���:jU�{y�����*)��;8��_�Q�pH$�욺�e���Қ�g�� 3�RgD�X�.�r}<ޥّ_��0��s���w�Ҋ�QL��������MQq��͊O�Rؤw@����	�)���?S�� mb�w6������I���S�����Z�~X�s�"�yp
-nl�Q̄Ya�<8YX�+��D:�E��}7�D����j��{��.����qbN��@(�p�!���,��u�䮠'�JB7�B
���un�;@�^�DC�y��!aX(#�ɄiU��ڃ�?�p�l�bn0B���nC�bfE���f�<����� $���FyE�ܙ��/J�y{�w�x���]�GW���=
�aSBhmG`Ǵ��@pc�h������T�͊��,m�w��*O<Ψx�hP�y`��_L���5���>000[��|���g�5q����iAlX2x�����,ӫ���[wF&��F���M|�!:����Є��������䐪) ��зS���jZ�x�ݏ�P��>�����g�����m�� 1Kcv@��?u~�߄����D��c{9+Qx�1�B�z�7"����]"�>M+�M\��ښJ�oK�����������KwL&�`7n[�(���/�Q�GtW7M�깨�q�p����3������}�}�1��$������j���]�v�7���I4"ᆩ9�E�Z�3i�օnX�I*�����
f���_�<��j�>|�v�nǍ�>�|�a҆��K.b��u4UVr�!ns����vN��T����ڐ{Ü��"$V�^�����k��w�^p<���,.���gK��%psC$o�sr��	<I8e2�:bF��<���VAb�ݽ�=n�̼~��w{����H�X4�P�v�ɨT�1�PY�u��JI�9�W��C���/J��C�W�jz���eȢn�9�����;~����Ч+�N0?m�:5+>ɭχ)޼}����z�sf1^ϗ�u�@���F�)U}�p��}ۥ�Z���5��K*���㸄�)�zz����L��(��O�4��*���l��]�!�%�U/�����v�Jnmiot�y���"���:�8���x$���$v�P�ڡ���k��O�h�>���{�(�U'�>3���m$�:*��5�C����bOk�����J�Q���R�~p��[Q����!##����Pԥ7뺮?�v�@3�Xڒ9�d+ggW����\1@,��[8\���z9���l��E���㕏|[eK(��BhW�4�(t2	'�ROϤg���/㊈�OOr4&�YVZ�����NW?2N�5syy-WF!N#@\?���FEj��Y��j�誥2�&�c*�]��j�j�yX�3���r��w�s�x����H�D��H��� ,@�j�fgK����zH�VUx�!~B{5^�_%�I��
�DRԇfErBy%���֡�m�v�;�o�j~A���4�Q�3/�*qx�!)�'}��V?/����U�4���^I�S�Λ�y󖞕ԯ�2s�A���b�O��O��$A�oܿ3�GX��T�<�J����&���@3U�[
�S��D[�H��XrA��<��,�ij��X'��/�bͰ��A��mϓKi��ӫ�:��X��dh׉��Su �����J�"~�E��K1�`�,4!�i#���X++�~��LD�YU�Qc�.��/��wΌ�`f��fbbbk���]����f�pVڑ�Ae���Ҷh{>D��́C9
5�GHH�|��G��a�;SO�x��ٿ>|J�t������^���[�?�w��a�uJggf����C">���
�M'S���n�d*�{L�ZBM[����9:��)(Z���&�><R��FGِX�yM�J��(��vT����� ����k:*��#g%���?�8j��n	;;�˽V��ڶ�� �����ڭ`321ӏ��D涋a�;�65�xC�򟗖����4�yJK�tJD ���0�A� |��F���Qr|�ome,c��z��K��O}mL����jJ*�)�=�6��f���
e���� ��Tp��H�M��85�G�X�#��g��NY/��1QS��`�;�7��Z�ag��5��-˴��V��fP�ɦ�vA��mk�Ą�q𫺰���&$�+��a�ͪ��q|aa>5���	 ,g`@����޼������(�=I��|�O�*���,��A/-�-���q�y��̥BPP_"�����.�MJ�O��i�*:Z77!o�k�@D�A0��w��{/�AU���������Z0K�i��D j|9^���!<�I�L�[��/�M�@6����hP�px�;|<�V3/Q���^���Fm=��mb!�Y��J=��w��X��/�Ә=@y`ˇ�û2���࿽�3+��:k��9<�w������r�2P_"Zw����?���9O~�+ ���w�F*6����aM�z���D��_�=s��%ʉHUWoŚ��$(q�|�#\ܷ̄�y�"Ž��ׅ���x���o�%�閊�H����+PQ�����EAcNsn��AD1�X,����{u���s�?�y�������.5g^�;�4�ذٖ���Q����BkD�e��-cO�/冠9������B���1���m6��lR8���<������� 9Vd�HqVà�!����K�r3�#�>�}csi�e�в��h1�N6i/�qq����I��j���p�S���3��%��2)�q�.�4��F٥���I^��o�K@D�O���N��d&{�IaL���zƑ�r��Z����(Fe=��-c�G���ex�sc�5���{�c�jtSn��.��)��jX��U8�1 c#2G5˃�a������~��#� >{g;{geA��H��S�y�u����H9c��-�(R��TD�WC���d��c�C��V�6d~U[����7tpd?>h����n��,:v6�ŘA;�h�Rr�1��LOa�L����c�h[��(6��C�����j����u�`��?D/?x�����md���❶����������}�`�Z��ç��.�N~
�J�Ÿ�Zl=�ӊ�e�c����9����#jhl,�d���QuOf,�Jp��R��3���&��aC�KP���d�+�&�Gyi��_Ph��:ޫ���;�!$q�?~#�z��w���iE�;9Ij�."���x�dcB��3)������+̌O�y�ih��Y})&+C��	���g�����r�p�6����B1�ˤEZ�5����CN�.I֓�	����..�%��3�zP�<�\�w�DWo�hc��*y��K�^n���O�^�])���s~���e�k�b�+C鏀׿�I�t�_|�K���eX��L�bb }�@}Iuyr��MӪk�ԉ88i����z~��f3E�xO��ۛ�X�5l�wH�NZ�10�F��һp��,;�#�ϗq�щ�
t�h���s�2�+�����$Mr��z�*UD	������p"t`�B��`ƏH�S���0��׻Z�(�H�^��,ĵӆݞ_�������T'"nhl�M꟠jm���������lx�U��/
�;4���u�J�^�����ݜ����q*���1-�U*���\A����4T���~�Yݛ�(8���R ����捸U��@�C)mg�X心��i��m"oBklf�����L؈� GΌ�<�B�2�M��f]K�Og�U��d&�E��/+�ʅ�V:�G2j
���:�a�T��PY��V���b�P��P�Oz�����Pz�0��||ϊg��kl�)��B�״H�s,7�,��"C9q�I!�z�N�@2����7���?���D3�����8�.��� ��U�t�~����xK�]_�T�3��m7<���u:�MR���t�i�n���0�8+�hK���2RZݶG �qL5ה�u�� ���#c_�]�j:Y���u?�gV�����5o�����z~4��8����m(%c�)�06n�n�W��;�����x�cK��]���N���=r8��؎eV���ơ*-��yx�gc�h9i+�p�DM��oa���i9W]�K��V؞����ܖ0����$�@rt�����tܘ�q��R��>��鿂^���P�,7h��@�.��1Wj㓢1�0R-�)9z2<�R��HuN�H���-��Dw����L�,*�����qt�wqJ�=��\�3�0���ڕ�81u>=�I������1�/�O���C#*����^>�n3�Fs��+��m���y@���_v��c���'N�� B����%��}o��/jߦ�hoH��پ��[>��m#����NM�����n�.NUo͗�l1�u��K�p{z&���߽���Ь�9,� 3�BJV����v^Hhvfu<?(�v{JNC{�흍��M��^  75bQ�q�=c+��{gw���
b�d�q���^e�oUo�:����t�C�b@��Xԃ�<�r�5V��9���E����V��f1��όO�9i�+^t��ɖAD�~��NM�U��]���:�r�-ץ�iF�uS~�Ñ{y9p��0�1->w���8̒cgvi8ޛ&(T�Ν"L�y��􄙝;kp,�P�y@������퍇8���x74gm������'R�|I�J[��`*[����\�C�C��@l�L�Q��Ծm�U

acMykC2ă�$����_���xP�r���(wD,O�������2;`��/��%�c]������W�����[B���,�ޱ��B�[g-��v�/��IEZs���[�E):���y�-4�!3u�nHŰ���/�[�+�"�o�R�J^��Q�\��E�J�M���Z�}|��~O�*��V�!R~���|��̽b��7Hx�����)���L���#�	k��*.��� A��xiOH/���ǧT+&�����4ĭ��u�������L�G@W|Ww�^��ޚa��@9���%Ϗ������� ��y��`�'�xBi�+"z�Ϻy���G8f���'�7�H����\���Bį^�4�Gr�G�]��bo0��)�����r������a&�	�3�v����֭�%��M����*|*Y\�l��$���b(>~����H��N5 @l,�\�n�˫��?�얋�"w�����i\��<�e"�˟��/��-T�]���jw��x���?�7�OSKor<�#9��ߺT
��8� �;������o�j�rMd5�F��(�ҡ6)��S���>���vswWMI���yr�7*�4,�7�S�iX��l� �|j��P�V�A�߿q��������'��}ݛ�Q	��u�t� ��\j<d�hb��[X剎�Z��547{BԚ��$�!�>�|�xg���+3/��1�(��-j�i�Ag9���}*�DE�����y*N2�1ޞ� 5��F���쐡\Wf��ܟY�ܖC	[N�d�{���l?f�d���
��o�.o����d�<<�/	��5Mt�9cޤ�{��Kt��"�t���)���rm���z�sf��5!��w���fF�^VD�{U%|$��̡{��:J�9�-�ݒ}8g�C�M/"bh�=�0��3c���*���c'���/���ʚ��1>?�z )�^L,~>��f<[f輸�%���j��4�9+��gdt$O�$����;rξZ����'��X3aV�7�+�Zl��qu1�����G'X*�|�1ZiX�oj��)�^���56>��ϟ��K�rd��H���tT8k+G�����A�N�W �O�$�M����� �g�g%E�	g5n�.����j�1�X/<�kCN�::�4���l�H�������Br�5��Ƙ��(pVx���f��������7��\��^�<<�� Dqpp889�I�d*�nTH��6��rwWi���q>c�F��J���A�x1"��׿k�
���YT�sN>juT����	3T���"�bT�k��%�������nlC��o����g3��i7����Q,Z`SL0�nh��8��WXKh����T�<c��S��́��'�"z���X�9N.��x]�O���-Q e���)�g}��g�X�Fv��-�r�2F������R�"�Tb���e��Pt��sw[u-���g!W�-�ӻWc7�a!��A&���c������<*����N5t4Yӳ�WJ6]띚N�����L�rK�~!ō#�exMQ��#�iD��c�%������-A���#�:'��rpt�'��}%҂*��������e�(�T�Ĕ�1�8F� P��'l@��F�M.^e�	{Dl�����A��J��>�mt����L�tR��L�jdj�&t�=T
Z
�?|���)Cۗ5�`52 I�RVS�F ��Çζ�#�Jr���S,��!�[�-w���,�Mk}l�)�G~�{?ҷ�EEE�;�ɛ'�}Z%t��[I1 	E|�I��|"��ߧ�e�e��(Q������=ܬ�2C_�/W�=.>����'�n�42�R��fa�����}��#&��sC���>wM�����&��z��A��5���1�;;I	)"p����YZ���I4e�K^��� 0>��O�������	op�mo�5fy���'bh�ci1�^�:_R�v'����q�$;����ז��פ?y+�����-	���ᇧ�x�$���yN�&l .@�!~�B�CdT������.�ৰ�R���*�b�"fdd�٥9|�n	�"Xe>�H������+)�m���W�����6gwvv�M�g��O���0��	����+jj��npϕNy�>���ּ'���XC�n���M̓�Ӫjh2w�Sp��u6������C�˼Z-�9F
Խj������[P@#��G�g+���̂N>��;�!��q��{8Ů�P�JEA���� p�j_�,�Ҽ��~Dڵ:���75]w�o�͚�q	8�������[�� �? �m�q�{c��w��ڳV.I�GNV[�)�,?��]����E&!�,����U��e���S���(u.��n�홏k]��D�Ʋ����xY���ДR9��Q�ӱ�R���ux�=�G�"C�{߆����}/�FĪz�/�LF�Hڼm^��~��v�k�6p��n�p�*㭆=%q����!�1P&�t�w��K��B�Hy|OK��i�)�2��8ژr��fKw������_M`��I�}���ȕ%:_�~��:�bxљR�&�¥{N��rG뿝��4$�ʚYhBZRNr��b��&f�֫��!C`prU���Xֶ_����Deʜ�]��#�r�q����)��9�N�3d�;:&%$��+�;ￆø�E�Q�������]���'"�W&�s��߹���y���1��:;��;(���!N�@�G��1+�C��_�C�k�� N�,R!�d��i��^����l�/�Y���u^
jt��F�h�K*&S����?y���y>
���.���=�^���0��|G>\O�_�_�x,�Ə������������t�qX ����4]���g��6���5x|b��ݨ!ftZo�@�[yE�����k�k�XX�w[���z�?V�½7�B����)�N����}��"�_�h���5r��wg����X8[��84S�d:2�׺��*>≯��a4��7<�]��}������ɕ�}މ5�jÅ�W{=4����j������<Nȹ"��p�啷w�����".���*�-�~]UU�sziM�o�Z��c�U\\�$h�>�>�eP�f^��۔�3]
d8�|$�"69�{�vj�~:�IY}k Rxb>�C�⑕a��~���\�� ]X/ѻ|�}���O*-	�����<�&O��� x8yu��,�i#W��2�L5������`x@>qw�<�X<6O6��(�f�W��/4'~҉�E&�WVbz̨o��R���8`v�tis8H�X1p�&^$(�+D�b~J���9;��q�Sj�x�%�m�"o�8�\��fV��i�w9�����j�=Kk~��6d��y�Fȅr��ߟ;��XJJj���CYڟ?o1.M��ͧ��2���8@�~�L.�Ӿ���#����(L3qu�NcQ�g�Mݕ���˴aiMM���k�R�ב$)�a� �%�ֶ�jy���(/d,� %�׺/���R��Q�l'�����S���,\��6�q��>��Ty��hi�#�����Z����hd��H˾�����Dٔf%�%��~�8qy��g�<��`dl������1�x���8�ů�_q8.+���^c�@�S$.9�?p͛�~�g�����z�L���ۇ`QQ�ӻ��=�&g�ť9���j��l����q�,��������-Ŋk�������ww����V
w(����0�3؛�����L����IV���ٓ�չֲi�)� �>����h��Q���ᑘ��sG��US�˝tJ�e����W�4�����x�����dz��@�/ ���A����J��5�����ߤ�͜C�q���P����ڽ��|��
��w�p㞔3׀��5�꽶A�H��\�Ws��F�����XV���PB�;�:�<=-{e��H�q|#�b�<'���=�U,zC�����\�B���aHA� �q���7�� �2;�xM�l{eW�Ր�P��Mײq�C!T��0��PqpDdǠ���*�.̭��&ƴ��$@�A]��"�yRQA���3���Ts�!k�#T�Mk�İs�����BG��O�{;F��B��)O�Z)Z$�*\�<`�΃NI�.���_f�t�F��7�e���8N���΃��au��2�(zc�GS��n�0�1�E��W��8�d��V���[ww7}��e@-tC�����h�F�ӗ@��+�Q]��%���X��Ӣ�>p��K��`,�1�q�b��"mHh5O��o�+��.Tk�%@���Q:�PV��f�+c�_�X;�OO$:�u'f
�.��F�ȅ8rx���$HIN����yw?b��)W-A]�0G t�=��hp��������c�[Ў�.���j��Ȩ9h�9��ł�aEX9HH����np�c�����l���$��yfkc�c�:�× @v�ɋW��BC����nq�^�����Oͅ����o,d��h��$��Z`x	x�U�~ ��^_�W�&����<7e��Hށ@�}����#ӧ�%�C�!�z2��4��T�a���B������A�F�᣻����sJO>�w�1���ko�\��{�����>�F�SrŮ~��>*"�����Z��i˂���񨂓���{b&><%���-������D�!7XGp��a�E���7O��K�Av��2�����guv�t���6�J.��Э��þl~��t�9�Q*�\;�#x=.23��'7�Q���'�rſh�V����	������:��G��NM�@/�N{'�ٸ*cK]O�r�L&��+B_���G���O���u���'�$g��&�Q�<����C���k5�b�O�^��L�[�m�`Wھ��1��}bL�˜�C�5T��H�#j�2@ \��s�  �Ƕ\ hȾ�_QU�G}��N��k,h=O`0�/䑙>,)��M�e�vpx��w����ht�P
;c#�\7u��}�f� �����I?�f��5��|������W]ǀFS!Y�5�R���`+VOfh�E��	�*���?�25�����Un��\���%�O	D�aBNNNY[G����=���y�@I���O衑�)��V����J4���$@4��gE/���9Ka��Ņ><�R]Yu^;r��zi[;2���b��K�ߨ#��O��Y]�M��������<�NWm���	2�g�M^�`� ?��_Qj+��tz��})���#�q��7;���T��z�ޯ��/�o�`=M7ך�||n_��h����� �����о}J�1;�~���{�����X��s�����N~��nx���!&"����CEµ�N:��r�W�����a��'
:��ba�m���l3��&qmy��9��h�ǆ�z�Yd}.;��8"FG,���tm��:�HZ��.Me]�� T�Q�]��~YM��|��|::ڏG�,�nwm��,�o����f��6=?���6v �'� ՟>Y[�����<ߝ���"<WI��\��+i8�`���+��:g��-��y�!��3��\�\��ds�u�cr8}�}S0]����'~���H��=n�����i�p�\�h��dW��]0l��Mn<�v�0�hX�}�}�@����_���<p,����M�ͭ���k��7��)�]A��o�{M7;K�I6��[ �vI��s�'v"�%��*�/8n��>ŗ�DEI��;MA�/�� aecԔ
�#X��ÿ.͖r^������䌜�|�x/#F�� f{����wss���>s.�Ӿ��Nm��.��l�E�!
�x-��n�!s�|��s�X6�̗���cT~h�����^(\�
�V흶�@$jxy��l�f7O���M)E봝�6-P�! -���+�Ϸ��mr:X�������K)ˑ�T� ��F��]/��<Ő��&�b`˶D۞���@�ݾ�fpP7d�է���[�4䅽}�<�,G��?�Akh54@X�)�ة��+a~�R�;r=�qqS[�莲��(��;��O��e ���I*K	%C�o�6�#��'y������zN~���;�K�aD�,�h�wl��B��t�����B�غ?�5}�j1�u9�P�]?xu�Q�[1�e��81��[�֡�� R[Ua(dh��72��;��
b�oMZ�AK���z��@rqQ�򻬛���CZr-�s�mUS۷�� �"r晵'�Z��;�E��֢��~c�T$b�1����
l^&4�$�3:z�V�3ªы��3�>'/�Cz5E�uY�
YҙЩ	���#<��{���u��[9���T�J�~�+�~]6��(�{���D��PxxC�S��+c\��^��G(,�y��+v__�ǧ;�� ev	�E����.����s~}^�J�1w;'Ĕwª��+��/i��ta�%$~��*W��'�o���𸹷�?��^l3׀]P��gA &_Y��;9r��v*�ѭ�Y��E�9%�����$/�f_j����ݟWWOW�����2��q��v�������q��!m���~Y1q���"x5`���\�e����*�tơ�@FS6�fzw��%��M�a�U�\1�,��Mt�LWѮ��Ҫ����g��x�O����;�}7��8_mO�]��pܞ:��٤�ku !#)�B����}�[ݚ*G"b�]�Ǥ���n���FM���iNN\	"����I��ء�x�2U	�u_?k�t����t;����-iK�r�ٚ�~K���N�4&Ua�����·!/����� ΀{�i�;~�z��^y�����*z��zH��}��S((��a`]���E�1`Q+ԝ�:xs}��/A���Tt�z������8E�(�әԁ0��?�3`L�Z[��� �u{�u\k�M�zy��r��b������-Քtv���0�P@{�9��Y�����������K�(=�9/�D(���u���۳�f�;�Eh���&����Ɵ;���:������?z��-��=i�Q��M��j#��x	}�ᆩb�������_�Wxq	��ߏ�ʰ?�uo1�p]o{��9�ω��I��:SXG7c��;Z����P[>wH������ʿ�~5L�/�]���/�j9B\����[��-8�JF�a�ʹ#�O[�}` N���6/;?t^12"���6&��q����4��Şo����1��	���Wa�nt
�#[G���j
ǋ���ff�Rxp(H�B��3�����u�6g�=����&����b{��ͻ��f0����94}�	�x4a�OBm�eО�W�k�De��U�G^�策�t��G5����i<A���\�UR͞G����cz��{ү-/PJ�\�īz:Bz�^��n��Xl��?N�����n�B�����_0�����{ӗ�c=�"�Pw�
�V�_.��ޯ�+�:��2n�:�O^}Vz=�hÅ��̱��L	� Eῷ�2�t�]"���m�qdB�'�wI�c���c[���
*-K�j��~���:��E��N��l@��APp�"jj�02�4��,���|�E�U���ܺÖ�+�lw�fv���/oTdT�ɝ������H��cW�y�U�K�~yA��/����A�b�ߛ�O�6������u�Ȇ���fb	�E��-�X-5⨋ߊC> i�`RV�O�g�{�|����8Y?-���t�m��������t��}r���I�o������3RQ�a��<7%�Ĺ�[L��G2�KD����>6��T{~�՚~�yW6�b��K�R��`cN,�d$���֠��-+�k���l�!3�nz����}1~����ނMO��W,&+���>�u�1�������9��5����C�
����9�������6Y���C�|k����N٤Ҩy[���8������DA���uzQ���N�����.�K%��'��@�%��^�� ˚��^#˽�J��\���+,�@�* ��+���kB�:4�z��0q	�Y�d*��I�-R��B�=!�����誙�V8)s�;(\���=�����h�h2V�_3��HX�P��ĥ����f9�[jU)���q&S�c2{�i���Vd0�8�:�tw�vuw�EE�.�I��+�u{j��H�������X�D*e����n�¹��$�O ���Y�����u�B��AռN����t��SW���8+'�/��z+�F��R��$F�U���{2X�y��䵧�]��&�4a��6ܞ~~���?�f���������@h�K2H�4<�K���/�͚״�*��ؿ��gegMak���gEIϚ�%O漆X������? -M�Hs2����H�B��@æ��Ec��]���.�T+H@��H�ϒ׶ �����}��zs{�sn�/1$����,�ןWF���rV�n�#.��O�i���B���$���#�( rm2n%�O��݇�p+�T>W��w<�����aaq��dl���� �:5\!�pk���֫R�Qj��5�,��:��<���׺=�'��g
�%��/���pa�7���b����I�q�)q��k��p����I�N�tr��3�kaг��2[c�R`Ķ(�SAU�Ċ�Q-j::i:���HH��h�E���E���N���Ra������i��4�կ��L�܀HA3�
�ة��2H�����S^݈!�̜-O�&�ay�-�~�I��OVz�`g��@��s��Q[:��I�!�<CN<,��fq�uDY"c>p�`�Q�م�!���g�way)������L>�=
��8KБyf���r�vS����H��) �<V$v|<e�wW�F%��Q!�v�ycgMU����"�>~]8ݵ9�B%EE��77M�M̯c/��|ɀ��ּF�Q�#�|��'�,������6�i_��ޱ�C�|=�T4D~ʲr,6�?hS�Ҫ�V|5�E!(�lKOjzڟ�
N��o`R!f�J�|q��0��g��Ťc������yjg���jfa�l
�����$�:_�w��b_^v�ڶ<03g�uqih��:��8h5k�^�\rG�踉����J�B>S�!���Y���sL�&p�x�o1���Ȩ�Af�IJ�e�����eMM�4�j���:�Ξ��G�6K]���咬�D;�0�Ǔ��X\�.)�]�vG3}��c7EN�v����}���������ǽ**�]~�!Kn��/r�����%yl5	́��WeG��T�G���B��������1�xCF�oT�||ܾ�	�R	�'�%��-ٞ��9J 3�Y!l��i��gE����<��X)?�,K_@^wc�~��<�竝CZFb��0)Te�����|�W��L)T�S �����|
����E�$�ۂ���*��7%#�?y"P���J���\��>]�t���?�W��HfL�M[>�k�W�[C�?�[U�3�T���QѠ�<t h�xy����R�՗�=���i���%�%k BI]ʐ��J�=BsYY.#�N�L�(࿱{���z|�?-���b���cH���5��=&��7��iW���F�ʣ���@Nļ;��?�A�Fô�����n3|kk����XV�)����(9|%�H�����)W�mCZ�i��t�ҙ�񟪤K~��[��8p�lh�&)��r�3r���M��L��N ���h�UiV�;9��6�w�o2l�A�X��X=�Q;1B�P�������%:�o��[�Ād��0Qu���ecv�ه�ݣ#��p��Ń�67,~�r�:}N^-�wZy�d�=qC8��i�!�����f0��_DR��p���d������PM��YhA5��_����U��B ����`��T�$Fh���4*�v��f� `�..��4�����L���ЌP�JΞ9(;���V���U<.��3�ժʴ�#-5=unvv�#&��ᡂ������<�T	f�-#��PC<�󚺲�����7o�n׏�.����\���f�\��0����iA���Z��6����bz>����k�xW�f�O:[n	6�X��d=����9�҈%r.��z�	�j<������o*����3
C�f1�'ĝڿ�VZ*�`��V[����D<��zl #,=y���74Sm9�����=��xK�灤�L5��c�c5�=�����r��z������#I�<@��>6�^toNq�g��,W*�VG|�`��a"a�Y^��"B�{��'���,�%z��q'9#��J�������%g�2-�ώEŚf*�0��4��[(���GS�'��#,�T��r���M�������3�M�3�L�>�@��{Q�Jğ�0Q���1T����	ɨ��?U�'�V2��� �\(ň*X�K�.(��s�d�*i(��W��]����} �o�#�ZNb�IO�]zzj�����J��`��'4��3#��X�**��mi�z:���YS'�H��暈�:f�u
�����������#	G��Hp22������=P���d|�yx44X�i�-�U�3Y��u��C��F~����#S̙���*yx$�d�u)r ���p9���X�cc�^)�i��v.�> lJ2�¨�he�V�)��ǻK/�qt��99́�(�*,���-�����䱽�Ga��.������?��Q1�1�)C���!LL>*�i�)S&��Tlg���ՏA����C�m�/��K���+��1����H�=Ntƴ�Y=�Lή���%����4G��uD��9���U0տ�D�4�	�NZ@��+�N/���o����&�G�/�ί�$��5meڝ���;�㈌�VEV��h���!B�p��� ٲr%ǿ�5KF�	d8^�)P�tLJ{�b����(���X��?xa��jw)�/��e��e�U��%[A������CU�N�����՚��2_m��}�?t���	���G>`V߄4��mΖ9Y�H{��j��օ9Q2�[��7ڌ	^$8,�Ө�����1u����l`�M0�.�u�ðsg��g����)�졍an鳓L?�2��m��I&��Kb�6Ô�����*s	��T7^�S���T���l�o����HHZ:+eF�w+���;���IA�+�����z�r-]�/s'�#�!~r���wwI �d_NFB�|��zf��P���3ZGm��!��܌�'�w��@��o�����cr���J��-����88U?q�l�dj��M���� _PWU��~��ʪO������/��!/.^UM���������������㺒�4pͳ�g��N��2˳"���E��-_=���Ri) P%-��������C�e^|v��'����D�{c�ڭ%��<�x:�Z<�z���!-����0W6�I��1!�	��r��#��O�>,\
=������h#��S�D�5$�����c���:��r�GL�GTwJ��=�Ū�ݛ~m���y�@�z����f_�cwߖ@���S����ʽ��c�#o���>��t`@�A'�V���^]�ԑ�`�Wgrp��>��Mg]7�6�ӡ�2�^��~N�|��S�?���k�hTJ�4{_a��4�ٔ���Q�5~!٭6����
�����U�{�Q�ތ�ۏ�Q��4.S&stz��5���/Z�q5.�9�^�N�W�z �ny;��_�N�$��� �ۮtyߝ��j�c�8�#9ڝ��.�5~1�oL%c۽������W�#������	�ý�8`{qx�����ħG�A�?,���t\���OH�_f��8�
�?������y|�+��4�$�!����Mߜ��3*������w�H�Y��XfIã���X6��ꕒ�z[�ra_���P�#jjϑ�u��]�S��F��Լ��i�^���K�ji�΄�!�^eUm�bl���'�衒ꚬ�5��)}��]?�LD̂����ڒ��Z����6������%I:w*� �e�wd�n�>[�Jpa�T:%��ğtJH�<�tî@&K�ʺ�>74�J�����45*V��JɈ��
jY��>k���{{pJc�r'\g�'>RK�%e�F�}�γ*N���+�9s_�X�;!�F`�����O��{��]׳���qn�lTI���7#Y�8���ó��j[�������=��;�����=�wcc3=��-'5~��+>�~�Mbo��'���t��̄�k�+��?Š;t�ddeR��^6�na�J���لL�#�&�Yqw+B�ڝ��'��|���9��y�UE_U�$����6	�v�����,�+14�m ���URXx]�rv����RQy�8�D�YD;F{�x]\X�S� #bHH�G��������NO��[D����v�x�.ge�lOp��+ψ �4��� ��3�GC�od=�����$��w{��&&��GCO
�HT^�8���Qk騈��BRPP�bb'P{��Q��w>N^ǹO�!��Ռ}F����R[y�S��U��ПdD�ߓ�g�K޺�H��	��|�_����ov�wtv����
9���UBemmy]ݶ*�摹�ǿ��xy�����"JV�\2)��t,�qV]�h9)A"K�h�:�V-�����ʚ���ނ�Y|/����蘘��{��6�ĵ�����J��L����ӯ�Q�c�\�q�lm)hi��=�jz�G�qN�V��Z�y�A5�A�>�90��C�S�9��"�7��<���x��xA���{$59aLڃ���Hq9�4�U���Q#�^h
a����f���9����
Nw�3N�_��z��S�/�-�
f3��FX�ޗ����&�N�e��]��VP(+�;�q�lH�q�Ij[��œ�����m�I��p����KX�����P)kj�니@����񸎎O�0
��T��v��VV��0�,Tɧ�#�Q�%�p�o�Ӗ�gO�I�p뱰��'y�;�ƭ�i��(7(��'�8b�3�Ѿ��82�nz��Wȗ�Z��Z�d�YR6�S�ٚ}u:{Vq������g�Iq�o� H�~d#�$ը�cF#�?��6zc[� v���#e�1��ې��\)���t���L/�%������%���'��,��L�4	����U�K|S���=xƟ��L|r�k⪔���=�������X�A���ߺ�E�~m���҈ǧ�j�Y�Rg��V=:���k�Im!_ 9N1hj����Ņ���<���`����4�xeK��O�"j����ǹL!$�\e?�Фԫ�i�~]YOLK
﮶+�y8�+D���=x+��|:2��ut@�Y[S�{��e�W�1:E�\��H��������O���� ��W�����}��������b?���ȕ��G{�<UI�כJ�I��?�����n�#}�����g/6OXXB����l�`22m��l��6�z{)--u9�w�Ej8��~��â|K�������� q������W����Xiż��kM��,��d���`��Z��Ҫ.���R�M����M8l�n�v��~��
�|>���DDJ�[� �x"*�(����w�na^QJ�fI��(U�|���R��)(�~W�n�oL�.^c�/��1�y�}̊�r2��c2�{*mG	�/u��G�6!s���ν��\vE�]�XN;"2ƹ���ަZ�u9�G��c�=�����g��B���a�+��x��.����d^^����F�7)����_عy�����j�g��͞��5Z�9�,_�!�2�e������R�LK,�pK���ޱ1�a*
f��4�E�w�Fhʔ0�,��Ϝg���ODc����V��ӰFH��x�@W�Z&Y��\c�O�9���~~�����&����J�Jb���ዩ�;��*"���&b!l!"�]���jF��B�-{�k���|$Y�;l�q���tL��b5�@lau7r0�XG'g���|�!"����_��;8/g`�����Dv���f:�� jK��F]pp ��?��v3����:Oi�^ �x1$��^l4�&~��1�5&���~p�;�@�a*\W�Vo����$`؊���OUVhh�_y{�_������ͅE�s�������;����8�<h�h���X�C��9���=v ���}n��?��\maIC@0������MEgO��f,3��W��J��PT��MR��w!H��*%2*���3b���SWA�FD�����ܼ_�oJ��B^�.������!n'ј��c�	:�#�Z�$I�T>GduUu,:��7��F.���}TD����j??U{G6+s�7�bN�����㹦�x6�<iiC�tǻ�����iS�k�6�k�Q��T��]��#5��m��,���f�G%&*SR*�^Щ�/���MNA���]LʒO�p������b`J>�X�:�B�[FGFGSr�¤�	��޽�!��f�F���s����И[ ױ�������I����q����G�g|�:	�ݯo�~�=4ϒ���k��:�=�zF����@�j�>b�������P�V-ih�[�rS6 )T���,�K��P ����[2�||1ב�.l	.���9��ՑL)�k�$���4)��_�99�:g\"����*n������]Z: ��NLUWq"}{�_��w��P�*Mv�������լ��^Y�Cؽ%�aAyxh��š��K�o ���O�"���IY2x�V�$��p<���&����ȭ 'G���|N�fR���7�kC_t�Ե�aL=5ohs2��Q�PSRΕ��p
<�')���PJS2��Q�o��)��`K��-@�.�����6�Z�|}"����a�W��O�˛��3�w|8����7ʝ��{�7eĭd�ar�����x$����&i "w�ֵ�z�O��r��8������o�!�w;������F/t���þ4�3����=<�d#������tT�;���i�����ݩc�<�Wz=�q��5�rG��_�����v�&���Bt���D��%X�q>�FHx��RpI���.-aNA14t`AHA�2?�'��vb�@�'�"T/���=>�sF#���<:N�=Gu�E��r8�y�~v%�����,R���s���]�Б�;�5��~���Gq�7+d������%%��mk�����Nag��d��~���v���`p����m�Z��	������pv���!k1e�u�K�oVv��E��1�2f(Ҁ�*NT�P=����&0��#��9�B�`��ޖWT���*�2����5.RC6n�/��6�%ޞ��37|Z�jFK
�����7>#&؎x�xK����%ϋ�3}����\��N�ʪ�F9)15:�xs���(g8|����{��F�f��ނ�hxu٤�$��q��Ɯx/vO�S��\�Ű~�
�� ���WT�e宯��\:9�4��/F��eg�d*��KxFVN�8�7��4k�YY���=��$��5_���1��2��G7�b��.������ӏs[k�6Iō�{�[�> �7�w�l�X�,�RrW�H��B���7�dwV�`Y��W��UY������QbV��	��\~���8�M���'�6z�x�����jTڽ:��y���xF5��9ȝ�z�'�������θ�/m��*���H��U�%�=�JőK���D �v�r�wOz��P��{zqQV�7h�B�DŚ�O��EpE\]qD1�@]�P�>Z��6�tYM_;�b)&��0���v#��T��u���db^�dUJ�6��=����?�����Rd��Ťd+��~VF�[��$�67ؕ��31K@���d.v�/��ι���~��x=;����4RRRbD���^x��\Tvq��H ��B�F8���002�RS'�!a�
���6v����������G�d(�EX�#�j	,�eo��T����7�)oj�D�oǚG���L����XzE�kA�����P=Fws}S����
�$l�ȃ(�1J�@D�,JKa^���շ7ѥO�>*h�D�G\��;�B�]$ͅ����ؖ-�)�A~+q��g%���!����Ώk����I:�m�hbѳ���'1���n�wF����!�L�F*#c��e[^�3yh�^�ә8��{�B�Ǜw�����G��l�$riEJ�
nL�=����e+�s�� A�8\$f��U�l��4��zƤ�U�߷9+/�x�!�������͆���Kl��N��{�εS���1���Q���֏e�-��[>=[�����~�p��0����"}"���ߢpczZcJ"P�m��{�g��� yxx�: �tCu�"�E���H�xv�����3��:b2on��]��	>��+y�]��<��p:nGk봕���Q �f��P7a�|
EA��#�w�ҡb[��fk=�U�����f*iiI�x1			E[��wu}��#���!��߯������ ���$s�9�>�.�-iG:A;.-�L�n�LdC�%���ߜ}�ͬ�U�矟��{_z����RSsO�>s��a� ��K���e��>g=#Ն����)�ê�wq,�T��Ч�ق6*t4�b�ˡ��"�I����p��MI�[�s*&�jn��B�Ԃ-O�˭�/�O�o+,���2��s�f���I����|� �I��-m%�����G��I�4�>�w=�]���fR���fS�~��%����UV�V�7��\8u{;�y��͌�cw�����F�`�(-FF�L��:o���kM��8�4�;7#�������X�n�TU<�_o� ���ӫ���?\Ǧ�Qra���]]�O�z)�o�3���Fo-/he��8�T��<����Zϣ���2-��D�d��ك�OW�}Q��/���$V����}R��F�0KZْsQE�����Lٯ�=�����Jz>9;ٵ6�WL�wP�|A'���$��#Wo���  �\'�XF,�����1?����e��;]�j��<�{��+��QX�svie����wLVN:�?�)z:Gz9����	���w��i�����~�P+�3*�|p�.U�԰�=�n��f��ښ������`���jem_�ǈ��A�%�#*�֔�N]�޾H!穅�e`O�IJ�A�$]V!'%4~�pw瘷�h��*�M���Y�	���2ls
�q=
�l9�\$�,S�S+�X��Z�᦬0񡯤�(FG�<�i�V�r���ڣ�e��HM�b�,,�DDBg��S��~_Y�h�X+<,�8�*k��*ZG(�7�tg}^�@̞}����_��w������\�O��Z�Y����������Hط���ZF�J���Ɲ}�!	&��e
���p�!�k�t൩�є��o}U��|9>�5�dH� ����xw̄��)/>��������n㹶s篡�o��V�7�'JZ�|q� ��ư�a#���]�Z�m�
������'槝��U8[�z���U��Ϗ���}Y�;��ַ�;	i0o���L���w� y)�Lq��o[GǑ���0��K�B*J�(�}�f��p�c�o�b�v��l��Qj��{ܘ��YoH��nކWR�X��,�lJM�1x���9�5v��|���be��Q]�ۈ�-!�d�r	X�OP�	��YXB�Ų�W'�nrք��P�Ja������,*q��Ҁ���e�*��w-��--w_9<�M^J#�����R��{{���R����"$�	ͨ�e��}$h�.qq��I�n��,� ���� au��III�Hg@+�*Mf�1L�;����,<6���1�O������%�����>����ϊ�����F�����q�7E	�P�>�Qw�d-U�n�A�6̍'K(V��d�fƝ�0�BLd�F�2�}L7��=;:�ɦ�ΜL��h0��'�&O4i��
f"+���ke�Z�H��#"�{�B����X#���Y�X��S��
�6�c�0�4çڼbY[�	K�^��܂��_�f� `[YMLz�0���~��V�'V���?����z`�#���������:ֳg��W�m!+�i�9Y�u�׃W�$�x;���z
NfM�ܸ`�	^S#bK�d�����,?������B�F���4G�ಟ�K[4�s��}C����y�9I�.��Ґ������/%�߱����lP�"^^�NT�D��0AY�}za54�,�˻v����(� bbJDtk�o�\@CE� %�= +�����gVX҈��e�{	�3�bԛ,�%ŷ�\�]���S�'4?~��/T�q��5νY��j�6�����Z�@;���h��.\^ʵD�Ӡ&Ϊِz��)��z�;h��L�py]�>�
�"�_��.]+�W6-U{|��_W7�����>ǉ˸��S����I�R3LDHaӤ��ZIJ��r\�r!�I�]qmyv�	7l�n�x˰�[�X�0��2J؇�g�A ��-��_c��u6~w�%QWV"��]6�����r��I4TÛ��P=��_�:\�J��?Djk�fƙ�4���T���0$�Q���o�@Hq�����v9�-K�؋��x�O�P�^O'�|��-��b�N+l�,��Cg��`Y��>&q�M������~��r���hs��/�H��_]��������9/?���j�?x�R�"<������n��"�|��^��g9�Ac��xw���a�M����i�~Q�hV��s*=��>�U�6>�x�Ǒ����@���"���)���O�� �s[�|��i����O�Ȑ~�sO�Kh���U;Q2+��b�`3Vb��+Za��T?��%���@�����5�RP�����O]G��v�ش�Fy�X}�J7����j�Y���*B�Yuge��Φ�'4"���q���M�m�}G���Z�!�!����0����!�N�7x�rJ�?�J�O'�ZF}����!Bז��+Q{���W��c z��@g4�tD� �yo|r�C&�X�L���W+���g&�<�-��]��(9�Q�d�Ft�q�n�=k9�N�f+��U�k���2u3\k^���?Y�XDy�-g\f\(!�Ip@�k�v3z#ŝ^4D�aE�k��.>_ֹ�(b�]˕8Of�=ٰ�E�mq�$�/ �M��N��}Ɲ�Raf��@B��1���!���rLY(�ܶ�@����}f�eR�(B�ٿB���&��'�����K�ٟ��� ���� L��e񅨧o��n�r�B:O��q��F,ۏ�XgW�o�V՛4 (��ޗa�ȯ�\�H�eE�J���e��d�Z+`�kL�zق�~�,u�§̆���/�nm�(h�XX����Bڰ�Q���!�mg��8�Z0��2lF�7���*��BAe��| �����'>���ʨ�Z�R��!��>�0�)(�_�M��>�C�ٺc���-nܯ�c,�ư�03���a�-�}�������?��c��X7E���Z�
��������ܨ�!��Ƈz�.E�Ȟ�H"�U�G��2��u@�\tm}2F�zlD��$���+�I�z����s����!0����u�J�hA��\�x� LC2y���L��}���u�l�P���f1�8�����]���i�z~w�b<$\��e�J�pxSL��τdW��~���)1		F�.� ���/N�dK��l�9�'f��~����)�nd�y�Mxb���<\��9A�{��Z�mrQ��9��*/���kvy9���HK>�?dh��YWN,D��Ą	�rW��1DB�]�d��7K6ҳ�+���:�����ƕ��ZL!�r$|�N�`{`rppIMWWVJV&
���OUx,w�r�{�<��L8��y�"�!��h�0��.~uF�[�U�xfw�>d�L1�����:l�Z�NQi���*(
���~CI0[Ej�>�=~в��/���K�e�3���]*�Ӄsrpk�BGO��K�L�oUkPl�`���`$���Ј��C��V�^:��Qő�r�!���n��2�)pe�p�������-z��I�P!�{ 4wop@V:�s��w�7V�Q�bbZq�F���t��oȢ5���B8t
"ɳP%��F�����V�_�/�I�9��i�2O��V}�3���B�`Y�p�l���IWG�v��X���eq��kqwww/N�b������n�e�.�����s�̜��'�ϽI&���<ȡ�c�����u��Vlx9dwm#(�L����$&F�8�XiБ	ql]����JHI%��%���5��������0@���ߞ��B�ww�\�F3���B?��*	ll�((P��1��lyr]b?i���S<�9�+ ��*N�^[_�n�'��y,U��V�\�e�&IM��ϟ��]y�&gټK�sK������HhhB&ħ��7���]��rf�n�7��1HX4XX�JZ�������Y��a�O$$��퉠���B�3�:����cm�����f����U�wڬڞs�x&c�w�{��ʬu{�����+���Z���<h�0*s��q��e1A=WȠ�3/��h���_)0UT��zz�����Oe.��j���\��HG��[�{���R��#v}���wwMU��ߑ��u#�P�(�����v�f�y�X�iŉ[Z�[RMH�Ƣ-��[�^��K�� ���S�פ�"ĕV�c�O�����ݺ�C���?~ILLW�ڸ�m��\�S&E���B���*�����Kp�*��U�|�o�a��c�9.���hr���h���D���h��<��j:'cp�w,��ɲb��0񿄋a�@N[��aE�N���?�� �G#%%��ݕ���6�Ƌ�lr����U��;�<#8����;׶�_،s�ەU�>lPaq�֤�F1%�RJ���}d�R8���-k��-�O�(����H�ʱ��T�:}�3�$�9�AkBfqb�#�����\k*����;��7���L'355�����a�[�r�P���$���3ѹ��#�V��1�9�J�S�D�z� ��������UL�Gu�1���n���F�!P�^�,t)��O�RRR�r�`a���R�[?ȕ��5{�JQf�\�t ���7��>z��Ku�`��iRU���o���|����4k[���l�V�|=�@�Q��?�'�}�jh7��ni�-��ɍ��ך[q���\_cU��!��K49�H�Ə�W!"����sE��^R0_:U%& /6��7R������7Wicg�B� �sS��A��L���=Wȯ6��Ͽ٪E\��j]g�/�p��ь�`���=5������P�ڞǉ�Y��5���w�Ë>��w�T49�󆓒f�Z?0��ީ���+�.��>�C��G�9+P�1���N��͝�����+_T\�0w�t��E���:(�֠R��������X�5w[E\�Bc�+A^ҡ�N��P���B�ٔ#Q{<�Dtyy5��LyuX
'f��|�x�۰�Oa�����4
���x.�&���M�����3�s��)S�jZƬ?�ȴ�]���P�6�R��Uiy�!?9����+��<��&�:�ݟ@S��4i�Z�w+&��Wi��4Dw1]U��#g�����J�GE�S10����=����Y�^�8�;�2�
�AU��+Y\F~������J�ߩ����r�a�ἣc�p睗������f�;(�(�<�������|���{�%�����>q���k
�RPq��4����\�AB���X	&�t޼4`�`�!"���Ʌ@G��c>[�/���y�>􋰰�{{`�.�D�^�K�ZPYa=Q���;���� }F�'��7�>�7\/�x?{/��ˢ9�hP �:������m���X���u�8��YV��v�(��7K���u�$e޿?SW��7;������nl6��p><=��]o��)-G��$Q}�XX�{�Lgrg~Qa1�"	��c�Ȣ6���ZZ�|�D���,X���߹����QII)��n��T�m�#pq�H�e�oϵ{v�Z>h�Jը�Ui	ivh�X+\���q��V������(����ƃ�f��:��:�}l0>��&��Ź{�c�<����+�(����4;�<MW�?�4��,^UA {���	�=3g��77�����%Tz�'�^!@ԊǛ%���
r�nnm�Q�t����}YCV�Xx�T�&$>kx��j}�d�-���vw��d���4iI���T{H�#6�xm���y������N:�r�=/�uu��٬�R�N����e/(�5P��߅ȯ9`rG<���^�cgg����e�F<�~�^��^�֜��2���r+�Ot��������wyyƐ|�
�����A�e���Z�2�^Qꒌ�l �|���lL|p�9��֋^"]�uL����|�/�/*��ñ ��d+�B��	w�ذ=Py�5W���\VJ=��,�IP�l�#���������~f�����c}�}0j��U�A��QD:��'U�:~ר�ϸ�3g��T*vK�����IQ�P7���.o��1��I��ٸ�b�����?�i7�=%�"��缻c^���=#��Ep�,!jT���,[��+�,���<1�M��������,����E��5W��D3�u(�AA��;�@����{TGՕ&,�����K`b�ZɄ����-��������%��2	W/)c#�.-Idi���6��U�R�q��n�>�����s�$�/�7��f~F��K�!������_�$��?�22ޓ�l����)�iu���}:s��͎[�y$��qBT��b��a�X�� m��<C]�[1i-܎�g����g.y@�W���^Q�(��HBYOO�a�e������ג������ύ����w�Ab��3XR�V�+�?���HXB%��&�G腕fo�eQ=�������h�vsr���T��<�چ��0����lm\P����dǚ� 3+���n��	&�F���u��Ȉ���W��܃�`��7
Y���+��ш��� ֻ��gk��j9Z�]۷e�����~b!!P�*��Q�:���/�6קv�;CZ8���Pߵ5]����u�}�J���g��YȈ1{����~�2�q��h��ͱ�Q���C"��Y�$`�	�[&�����^�klMKn.	''��a���$R�����[��oD	Q55����P}iy������C�P�YkNο����a� �4E;�툒����$#��C�f���v���צ����͝��i�7<��eQ��o˕�K�gdt<xU��9�F8M�C�E%�	܎�;�����0g���ŗ�A��&��$��ǔK��IbKG�]Ţm��(�3(��O��ߢ�o��F�.Mߪ(��!0ݢa!���PH��-AΠL'11Q�*�����e���!.s�H >��Ĥ�W5���gJ��n��Q��F��t�m����,'��o��v �	��.]["��Br�5WW��#��I
x7�KɅ�b�{���nH�n�������lK�g���}vv6�W�%�n� ��גԖh��^����F+��K��s���Z1>���l�X4$Я��U�L�Ig�S��ZZ�rW�^8D�c!#�qY2�E�~��C#�V;�0�UK9��<�\��E���P�I ��N�t�@��G���́�P�r�/��?ž=�㡌��o����Z��l���sFC�ׯ�QՎ��)>|9�w��=��VYU��6�x2�Th���⪿�!�R�G�n��<_��/[2z3TBE�1���Ǣ&(��ce��y�@MWO�{���OSlz�I�>�X*DV�t�?�|�Z�����A�bH w�����z�6��!@`�}�St�q[[�
-��ܜ�]Xwà���ͬ�{܇�P�!�D��ov��Vh�N���j����鋑���+�P��}r�R����[���1&"%�Z���(��[#�Ш˓)����bz}��������t����g.#7���%����wV�����5dvr��kv�ޔ��P`K6��i3M���x��#-S-w���{"5���{�8r9�%q��bi�yuqvf[6�4�s�����,���l��'�m� �B�+f�뭝%+	5�k����A�P�j`FV�A��l[8:.��x8K�X��t��9�կ�>m��v�0ۄ�ffE��s�9ט���)X�eQ��v���cΞ<e)(�Yto��]�q���[�̝N�K$����������T�qy~�r���E?��:wY2*r�.�"����}>aE��b�#\r�F �W�
���9$\����?��
�\l�'��Z�������ɼ>�X�)�豯I8�bi��5�Y�O���k������5~���퍶�Dg��?�<���D�r7C䳯�0�qsw[o:Đ�oʯe ���������lw?��O��k#�臛2aq��ˢ���	+����	�@w����;=��	#��Y���7��G����� �>֏fEf��F�u捤tڥC'�(-�ΨP�п�k���W�	�r��2.�*ݡ���ǎp����n��צ 3Wۤ�_��
,��v�����98���v_|?1�]��;�f~eԬ7�N��:�n��9h��	�ǋw���0	��C�t�����g�crP��7���^X��2���q�rE��0�Wt�cn�L��/�㓒��^h`�o���n����M?�i��ONr�>A}�i���$9���w:�tΌ��e�o�nEM֗�R�'�v�J^J�&+�������
�"o0�̭�f�r�?�		.��������w�V{��~�tH/��O�r�k�࠺|���@� [��g`���{��̙ "���ͬcKۿu��j�F�hoӲ���Ҍ(��c�F�	�N3auYGY�eØ�k=�;�m������4Dϱ5W�*����&���Z�cB�~�z;k����^z��z�������o��)��Q�#���B�a���A;�i��>Z�k��d�H�1����slO,���s�=3���I!�n����bec�GM�lsZ������ǻ��޶ɀ��N��$�f�C�����1�Cj̜�Y6�%8u���z'Q&��jC�Y��F@��2=�0#`��|ЅZ�
B!�F>��N-uz���%o��/�{�ղ�:hOɜ�1�#��Yx�9%9$�>�_7~f��Q:���`�{"�	&�����oY�9�-/o�4˱x�z{���e;r��bB����ڒ��\蝧U8u�1�~z��Qg�^���\_=ҵqܞ�z��W����uRa� �<O�w�?�0*Y��oO �Pn�%B	Ҍ��X��ݲQ�`��iiYK�}'�k��k�
BU���ș��ʟ�R��J��/߫s�46.^Mp�!^h{iÇ��a|������nbk����,�9#�(�?>��;J��K�4�����Awؔ��

����=3�X\<!&���&끮�L ��1��?��!���5����m�T�.��;cN�ʂ._}�����sK��u��n)�6��؅?��O��|�}�:�8�!
�d����8����)��Mf�d�>Vp�F�c�<3�բ�o�o��v��?�I��e��0w�8�ܢ�(+��\[2�?�v?�x��ܺ޺��ݩB`�p�@�j.SY��J���R�>qE Q~L.B���_�_o��
W��m�������_��B��o8f��[�F���u������{��j�+�/w��H�^^�lad�I-��l�^��o��[�?߁�	��T	;X�w~}��CU�;}��x�~�z>VR�ZL��=�o1�RR"5X���G7ug���f�H���̸�X��r����Tݡ]t���i�1�ЉH���>��Av���/w�hy��J�d��ו�m�_����U����@oo�A	:֙��:rqQz��>�[��h{EX��m��r���e�2�����?�x������g���yw��PPQ�k{`���O��8��&�X�5��ʲ'�q�z_��[_.Iߐ�o'F����h�\�5k,o�@Q9uI{^	{��ߠ �G����Gp�R���	��հ��el�_M9�v�wgY6����~=��,Հ���!��]�~x�][��xm��R*��0k�J= ~�h����|I�N4�G�D�v�$�ؓ5E�ً'ላ�lt(�xM���^�BP*Qg��1K�0�Hz�l�l�^�6f����0�M�	�j�`Ӳs(�ծ������ឥ�ҙ�(���.|H�����'��y�N�e�F��\MC�[�&��.�4�"����	胞�A�i�7���Uo�OK8�X��͈󤊦�׽��WzmFʧ�N�-����m�ָ.����*5�Z�h\��7ÒdCĒO?Y������o܎ޥa����j{��/�w`�|�mYS�rpp�&��m���@�B���u��3l-%�-`#�$���%h���*[O���9S��l�� �X���^Aj��ƞ5to���*>�k7E?GZ��C:R@��fY���G���x�hx��BQ�m^�D�+�R�d��_��L��(��?������R�d�ċWl�6��"�,{�g啭�#���Ej�J�w�k��f�eMjظ���"k��w�u��=���W�m(�t�M����r?�8�8/�nu�0��0&��õ���U��-2ִ�c����?��x�0b��V��l��tAs������I<a�Վ�����P�/�rRRJ.���j�4������,Bd�UB��w���3# �*YTc��v����!�������0@�ɞ4�$s�
ۖ���J�?���d#�4υ�{���&��׺�"o�l�?��+?7~R� +y�'W Ǯ�.�&�T�Kn�<J�VE4�3������Z�lR��@�?$7�R'k��c/�.��9��Q�MGm���Gs��B>��QS#��X�����G\�B�0Tk���/�H��k7f��!�'"������g�N��E�}0���y��^��{��/E%n�B��Aq����C-��3����	O�j���D��:b��^'�K�B��*)FX�)H@-�+����Zŵ*��S:Z��$rN�Mq)�h4m�"Q[����w#�T맵@b5�#���9�`��_��͊�#沱�6T6���ؒ�dq֓S*<���P.��1�,~��3�����؝`���#:ѡ���t�9�"3�ILOJV��� �v�~s��}^l�)��>;ب����7x͢-���s�'��[��_�8�R�0[@�։_����UD_�EiBr9���iW�Uiw$#����j��q����G��������<O׋�_� �;��L��]������P�Z\E�YΨB.�V���I�a|ۙƊ��A/���u�C뽷������8�BD�hp���Qka��܇��h���4j�U�T���8=����d(�����訨��_�)K�1�a'��굉CSd2i���&4#��
z���@hn�V۾�*۩�+͊�4���MğZ��M0&Yҫ�գ�vS�4�ʆ�+ 
h�8'f��>CiJ1�,�M�H�E� f���	�F{���uJ��0�ք�Y�,���o�8F���G��;M���7�ɯxQ�%ʖ�d9b��)��G:�Kb��Z��TKTʐ-�ɏE�o�tz����k��o9�fh"� =s1��)��X����0��fq-ēL��Sž�S�-2�Q�&yVH�I5Y� ����!K'�h��U�RQL�������R���h�Ek�� ra���ܟ�9�����Ў/�tF3
�֝@�P�;�EO	 �z�Z���Ԟ������ ��s��إ��F� E��X�#�BS. �� ��\��j���y�c\yS���&���6��I%��b?=+�M�yrc@���P�L<D��Q�hP�QԌ����YQ��8��9\�i��$��a�U�M"���4B.�/]��a�9�e:8|�Ժ��b9����u8�����[��yAG���|&d(ɜNLFַ߯C��e�AOH	x�3=GO��`��9����=��X�94�AVsw��~��본�R��*Cs���C���M��E�����g�]��mB|��h&ɨ��$L~0�p��d��-���F�>��� ��d��2� ���%��t�c�T�k��؄��B�u��]��aLNWM�+d����M���:�Q�����U�9�������t�U3��g��Sd1>���kJ,�pNH��h^��ggGW�t���Ўq��GG�l0���:��T�#7+��՗�����)L�c�ch�+&�k��L���������'s"�*o�g����^�)�L���b�\��z���q��QP!���d�#a)�9���f�o��g��8j�<�4Wɤ֎��E��	e��@��]��$#WH�?��9q�1 ���y�n�J֥���g��'DmboQ��Ɖ=:�<�m���l8�@�������t�*�%��ܕ���$���$�嗄 ����+ob��va oS�|��3C��O�p�m?%��
�����[7������g$F���ڔ���>�E��p�|�I���Z��i60O����SŎ�qaH���nы�Y`BX�6g�5�%�<E��3�J65;�El���RBR�CX/����-1g���	_;�zd��,.I?
��G>B�
�e���
��L`{�κ����dbe^ح�Ybnq�S����\��0��R�}Z�~�@�s)v=�"߹Rד]9߯�IU��^f�;B[5d�4��^��6V���2~QՕ�&�;K�n���-V]H�D10;�`jI5�{�*�PSvx~� /W�����O`X�Ǽ)�(B#Pu�t�O�P�Xt���h��I_�|<YW'���|����70��ru�;���;>>.X���o���Z�y]���7�QY���Lx�E������������LV����wMդ�`I<5���T����3tD3X�R*K$	��L�=��m��x���I�rϔTT|��<b��9�8�����H�:�m�+5���m��|�W8#�r	)LP(�&I����T!�o�3a����x԰?K��Rɫ�>��k����a�en�B��!ivH�T�X<"�FQ�Q����q����%�,�&۶&y����_d��%��N�?����y��V�#������+7h鱄��4
�����|�x(F�رlinf��L�T�4w�x��Mό͖��/�:�YHa��ux2v���e�M�D	�^:l|<ݟq�>_�9���32�0i^f��M�̜/1�e�<�xd/�8{~�0%Oe�M�\{a2r�KKא�9�ӂ����UAl��aX�׸���`��t�=�� I�0������j�
��u�f�<���5�4��kKNM+�B)l@3�d����/� �c<]p���o�m��ۼI�-�;���!���_��џ�nw��:����/JY3
gf繂������t�ޫȶ]]�*?F3�W}<��J�JG%T�S���b�[d9.O�!���Kb��_c$�z�׼�K��W���~�&�-�κ�U�K�tI�l�>��*���T*�������O��ڠ}du~�4H�bQp�nJix+��)�A{�s��,Yn1H}5Z�Z�Z6�)��7�봋W�U8����VSÔ2EQ��mБ��d���
]�	��C��;Vt���K��~>?(`B/�L,�xH�
DE��N>�J�&(��>����)վ��GYo�ǎ�|�:7�cemh}ʹk=}�Kp ݜ-��h;��r�d��"����y���ts{?oω8��,�d�������0qp�q��zWp� �Y*JT�!nWj��c�GNy00�i��k��>�������Ѹ�HN�=�=��;Yϱ;�.^&�_]�z�v���o�kJl��!��sj��&��=A?Z���e{����m�=��j�/�K'�ݕ��I��09��7����@oq�����M��3����(�r��ȑW��A-kB&��"t���p�n�5H��p��x��-ޤ*����%����8��K���ݨt�5�x��Q����}=ĥ��m7�1S:�u
��r_n��r��@������J��E���W�7�B#��~w�U)�K��^?e�f����<�w�������%Z��b+W,�\W6�\?��}��kO�"oz#�樭��o~�����hN�7:�Y̟�������n�ܶ�DaFзU�=�X�/`n�������w8	�'��nܗy�_�۶c�܉�sFH�bk�S*,��1���|C��o���jJ҈��v`�םs��o�0��6M�)r��W1w���l�����|��]�����bt��]p �f�;�I��RSg�p/��vrB������<(�Nə9�6z=��O/��À3��-9W.� �y�8�����!������A�Y� 0tw_
�c�~X�I,���.��ۯl �;�|U��Ty}����J}��_�K� 
zq����.��Ι���������5�Iw��Sǉ+�|����o�a,,ݤk�Ꚕ�K��s��� ��.^ӠD�`Q�E�Qzt*�"�٫רU�t���2�?#	�H/M]���E'�w�~�0$B���-?���ltȻДwU���<y!*����o�����vQ����?���� Q�F�\��{���wُ�=G[j�wa������G�)�2<"�Z(X��'���;.G�"[��vk^����Ө�eǣ&���@	���}�S�(��%�Zu�i/*N�d�l��c`ŐC4�)`�`�m녊��c1��d����r8�q{��g|�������upU�����s(+b�Y�q�' N���P"*N��7_�=󼥄�Z=A�1m�z�`�P�}�~Ds}/(���gw3eܢ����4���Jh��5��W�b��M��,�����^;3��w�޾΃��J*��R/�r!WϤ�p�=��/�#-׷5A�OV)����b��c��/����]{��iA�V��#�}+Gt@��ȷǄYb|yǷ9&��	�Җ�꘴B=1DԻ�x���*)l)��'��{����8�#|<�8�0z:l�כ��)���G_iN��Bj �n����? >�n�6��?1>n��l�C����R��@�6ҧ.PѦc���4���I��d�����R0��0����� �{����y��v��&�쳀O�.�#�їCT��-7n��]�v��'ƥJ��nRVV�ޯZ�Y�݁��`���C!u�N�-*b%s��W-eȟDK|/�>Z�E�L����f�a(����A[穃SQK������w����z�Uv�j�G�w������ΕnS���8?|��{�̆�o�J�� �_��@��łMFC���jyO�P�P�^���h��;��ӳ�k�\�B0y�'V��ͱ�vK����)��i=���B��V`��C���[Ȫ��,L�.SX���&���t9�����^c�@�x�����%�
6zC]��ڿry���d5�D�E�A���]�k�?_`"����'�y�ϰ;Č�����߭s��)1�RW���S�V��"C�ЎDTa�0��dô���6;o]c��fe�2��}��%�~\K�ȫO�m���6W`xz�q�NO�,�8	D�N#ޔ��6�,F�G��ܙv&�CFT⸛�����ǭ�S�a��}κ�oNNM���R&�����$�q��(�it D�=~���<�w�w%�h�B���z|�����p,�pn1v���@�'�wDj~�(Z��2"쿋���HG��g-B[n�I@5Xe��r����/�?�VIX�y.&���,��P<���*�mttq�5.�m?"2��v�/��_���_�v'��N� \�HDc �����eTȯ���Oۚ�QB���&�TN/;�9Q�;��&�j��Z��_N �p"r��)K�F	Մd
�88�N��+G$O��b�(9Zu��R���������p���4h#�������i�Ʀ�>7/�����Q<g)�j��Ru�F_��a@��荤�%�szn��ؼ	ِӣv����[��H�}�����Z���m�Q�y�f|ݶx�� !N���c�p`e�0"�!_%�L���X�)/I.�ῊjS{���E;r�9��F�!]�MQ%#��������Ց �e��v�J��`]#R됡��o����4ªx�S�K����w?��zyq�Ն̜�e6��������M��bG�z�iMuױi:�|,^*6U�4A�?�/�]���x���*�˓���� ��e��<�IO�H�6ck��T�'`*�8'J8Mp��mn0b���u9-�ir����'^��6��}��ƿ�|cٯ�C��hRg���n'x�<�T"~�֔�]_�RG�8�������#ز�w�潏�pp�'��H�\o��\������?^�گ���77�#e��?p��D�
�hv��r�����f��YYb�Z��G`8�����^�͖��]��d�]�k=��!���R�o��~�؇
�) ������	�5�C��r��_cJ��WD5�F{��	�߂b�o����kL���x�y}�1�����\j�O��7g���@���|�ۋ�W�Թ#\rd�֡�¶χgefkV�i)N�kH[
GuN	����T������.^}d��	&x�uQ�� �)�H���0(ԅ+�26F7}��dH�Y:[�K���}�����t`P�B 7̂r�|{��� #3S�U�4��hM��)����]�.8>k~s�K��u2��Պu��W"[�ҙ�۠�;�ם�Nt�Gr��x��k�
�sMT�k�X���E@�[�� ��18��`�����?k�M{�57I��O:p��>v���yİ�j;��Y@�㣎��*{��B�>�d���#.�c]��l��m��������Rü��_�d(Q(�������ZW$�����f�5��9�Ϝ1�4��Yʘ$�����ˬ�d�^�4�����G�7�g�MM���\�wګƗ5��S;P�E��Q�A]Y�(����
6~ni�0oC�	�P�$z 5+��R"�����M=v��{N�E�?�oCr��4c����ˮy�Z����v��"�i���<��Њ1;���M�D�\�*O@�f��{Xڥ%Ӱƙ8�����(�V�+��L�����<�މp˪�82{a��P�����
rl6�_v�Č`�?��iX�O��u�������-^���^�Р�ʦ:;F����R��<�y@��Jw���� �M��ul|��D�6�e:&R�����gI�0ɯ���'(4�)%�(�G�ih�E���(\�]���B�Y�qIp�P�Έd�,k�e[�r]]�5�.��C��mjq�y��\}�.Cb�=��~Ӎ�k�UP{.=��w�s��P	�*�~j�&X'���7���P>FO��u��{�!��gM��gq[Z�HmÕ�0�Y����\!k�5����~�P��Ttl}���^�W��A!��G<#0���g��^�z��"GD���I�*���
꺿Ω	¯�69��޺��?���nk�����(�{����o:6a��~gCW(5�p$�R���P�hu��ɱ�Ts�5~���X+���49e��D��w���!��k:�<n�i�ỉX��,I�l��)�����lD-���A���������b�١���_6���������k�0���} �F���O�4�o�=���Ɏ"�.v���E���RA^��~ӋeH5�	�TA @������eu�ը�,�f�4����𴋵98ߑ���u�~���8%�~>�𶎲`��Ûp�1W���ں/�����5��T�T��.� �K�F��\g�6��[�_��sn�a�����5;���mo�~�9y����ȕ��9���X֗,חZ��N�B�E2�Zqu}2��S�������:��T�w�Yr�����m��lH[w�J=;#0�suy5��F �ě����*(*�N(r��0�=�x��Imo��aF��SM^�zn��;�56_ �����&[�_R+���AS���6'��&����藤u�<q��wOȯ4;��j��6=�����v���@U�Hⱴ?�󓾻��!���ZD��uC��G,<��Nf�u�s7��aƖ�z�݉�}���
��~���WGb��� ������H�i�GV����_���S-����t�{��w'k���Q�	b��=}�^ɫo����F�G�h���������/ݩ�bx���L��8��SQ�vV�2�vE�������~��2Pɪ���j7�����R�c&Qޑn~/P�����<��5kC���1B�|s"IעM��O�)	���s"�#4�����s���Fyf����yז��)t�s�q����Y��ȁ��>��gB�{�9���؝q�Dj���,ğ�L�ߧ���95˔���CCsw��,��8�y����g�v��'倲`ni�K��Ki�D �1U�����sN��%�U�*�xfK��D5�I�,|�M��Ͼ('��.N{�޳�F}8�ϟ�a�J�S_��E�3ҳr,}-�#�~
�yL+�����S��
?�ŗW��y��
+4)�����[_\�g(㨊��R�T��M��>U@W�;]��U�V��Syn ���;/o
�y�zn�mRf�_��tt���ݼ�P$�8j��%WrL�w�=���ş�v�{8 �+	�r��{�WC���bS��[���%��R�m;����T�>X�����3��ީ�^Q���+�c�/���qM�/v43���E��PVjdD�'.T"n����?����&
WCL�p�F�7���U���,+�7�ے��H87�/�,O	�����*�D{�$�O��枾�;; �b<:|�uf@d�T�.�M!�*w���dEu0��3�n�z�� +6!?_wZQ�JcPp�����(%�^+�{t�A��m���Z+���Z�����PĚ���5?V�AeV��e���kQ�H�M�����kȬ����q,�+ԯv���Ζj�!H�w�G]��R���9�yJ�у1���������Xe���Q�Ɉ]�X�}����6����}��k�-���V����-�z����2�K�E�TN[3$��b�G��&�{�W<����7�X:u$��z>�9!r+q����O���G���=z21$����7��9��[t�2�a�`2����!&���2��+��L2YLw�y��� D�),�F�C�N��/��_B3��e���≽s�ۑ�YGU��>�İ���Ծ���8e�UO�B*���wy�F�&�A�̀�B6�?�v���RվÅEл�Exص��O �b,��=O�?�M	��f.ޠ�} 8��)JX�N��J�Mp�z��˻���]�a��g�ڰ�<��~�^"8��|z�i���+�P��U&U KW@y�e���3n�l#WM�=�H#��MKp*"8���P��g/a�$�0ֶ�RgH�r��&<|�A!5[V���Ѕ�M��}ۛ�+b�wT�Pd̦�<�fd:��E".PD�5o����5ո�U�L�F��kwe����L��掦u�P�=��E��K���y~���MD������PZ�6.K�+�6oAf&W=��$��"RX���~yY�h��+CY�?�]� 2��X1MT��О�go�D�D���(��������@s����@��9Pٜr���:�!���)��.O�EG�|{��GI��1���[x9�|K�wE���Wh��o+���dlpK(O@�]��˗���ug���Qew���j������N���y��.�^��r�1'�5��t�K�E=�~�<4є����Ӽ����~������vOAs@������h�W3���r=i�'��@�Y<��0���y2���1q��=~�N��$�s��#�A��H�)[��<�P��z��q��I[o�0���!R=��3�M�\[��^I�������d�߹����<}:��y/����vs��q�I�)�e������%�^m�,�B:�S?��H��e�L@�H����H��J�q��E(頛@��" �,�+;�tx����-#u�2���u^��E����a��8����m,'��P�]$�䘆z$-�P�s<F���Vct��������I5�(୆��w�H�Fs\E��A�c[ִ aԬ��~�����8K:�z*�Qd9끌d��~�%�
2�Q>o=A^rڀ��M��zz�K��	O�逩Oi$f�O~K.S��b[�x~X��o��Z:��-��Մ��L]��o��GH|�'�� P�@�gQ5�]��9���Ɠ��ع�\x����LYd�+-��5v�|�Quʺ��S"ʝ���2�J`7���4�4�_��E�,�\w8�m�5k�U�FhD�gj��Ǝ�U��{A�!�&v����*��Um�~y��r]I�<����<�9�T�TJJ�N�X����iec�W̞U�E��Yf�D��.]���GDo�����:N*r�����dqE��F}I�m!挖���_�9v�ѱ+���z�X��G��r�0liO��S/ZX�����7����vu9+����tু\����G#�Y�CTw��R��!�k��H	K�iV�hc�3�P�'�����B7�\yL#�"��Y���L�8Z����ʝ���NJZol�@��C�!��R���=F��%��~��cO2�]�E�D����x�2��"]�L�+t+��З�A�i�6#yN�����wt8"�+�F]:�L�'/�cː��]��3���|̒��y�[��5Ri�rJ�`���\��.��؏�+����Y;�Vc����W��΂7��W2m��Fe7�JP�R�g��g `C�W��N�d%y�6}Cm�O�]$�o���M�'��9ϖ��LD,�+e�c����`É��_2�6r g�z�6���]�;��z����	іI9>�ZP(���D����*P���,�P�cH���8)�jrt����>�썮B��>0(((Q[�g�w�u��K7�&��~�Py�q�8�x͡��,^���>��Qp��]M�f �. �5�iș�x����
(�D<H��L�}�j�J����9C%�6J��۞��	�ٶ�⺊�
\`�ϵM�q�e�[x`���{�%�E���K��宵��&�#h<`N�A���ĒB�ŭ�.��]��R�A���5���*mkyb˖֧�EY�l'�O��<�|Pf.��� [�}$���6�]>�ȌNu��j-��:�%Ui#\���[�+�2���s�mmb�Pt�T$7����|Y��P�(�>B:5*�gO#���<k��d[�h��>r�U�x�8�1$�X-��3FX��`?^����$����:@Y`�꾣��GJe3�6���v����X�7G��bV�N�b�k�i�?�^��;�@/
���((9����S�%+V
�2V��M�������:�/Rt
�u���Y`�>����ׄ�h�?%u�Ȯ$C��Py�$�>Fꚲ:�1��^��(=���=<T��ӷ�eVv�؉{cf��}��6�k��R!}lz��M��ʍ��o��>�I�����F��ڽ�L�5��v�LCUH21��������O��c!�,"M�.����';��ļ���L�*7�E>��	�VNٵ֟�I������h�/*	ֹ"�=C���� �ɟI+�����K��p2,Y��V'_|�����#����F�Gw�iFhA�~��S�wyB�������Ԅ��
8X\�t�����^�tT��h�)��3�+���D=�P�eA�
뤀+�¾����}e�JzUIE__�筜����7X��ʆk�(����kz�6\��'�I_�F�;Di,�<�F}�	�n0� $(�7D_7�����sE+�rs';&��?�2�x��&Z��а�nO�;�w��gf>3��;2n�6�p~��Hd+#<1<�;+Sx/�c^��,��ay��z�����{f.Y��_�X�8�:a�:9�1R��_������^��:�s��t0��w]Sа�/���#��%D�G����P�u����\rol~2�,�2���_��Bk�f F��"5�j�i�yUR^ݭ�̢��I�J���D;��؏�(�ؗ?�M$� ������
'��J��葏���cr���=fey.�G���Xρ�ݺ�,>��Ơy�(�,�>u%�g�)�	2m3�u�{��\FCΦ�8� ��ð�ҕ���<��>���`�?,�EC2�5�o=�����f��kxQ<���
Lui��&����HK)#-���ƌЅn��ѻ�!�ώ������/�^�X֎�޾���#����s�
řI�9�i]�H�/��I mn�O�%Esj���������d;��)�>{��9������u�vI��n
��������ۛ__�����a�W>\ش���dM}��]LU�W��Hj�a~A����ϴ���:ܻ���2

O����tڣ��%�d6��pu��LKG�d]���=����O:��>M�2�x�Ѷ�����b7����
e|�N�KU�3��>��LMK�O�g�|u�qWc�cz�9��E�\�b��v��+(K�d�x�[v'UҺɟ1,ç�bo����}1��ֈ����5�Ҙ#y0��O)��O���k�e����U��q�Mz���M2���eSf�}B�^%���(�[��`)��������و�yyu<�Dp����~��� ����X�/q���b�YHx����}��տ������I*X[RS�~�o�[�#T�< �{x�C�����>�W��B��å��_�}��>I�??m8��&��71��]\��f���񉓱c�cWl	x�+�7�ֺ��o���L�'��9�"��%ƛs6�����K򀝾EN��/�F�x�ݧ򇰫�b[��i���vҎ���ƫA7�H�Ɯ�X��W��ּ��/�RC'L��o���}�,�,`��n�>���/g��l��9D��*)�:o)cOM;v<��q�(]!��UBL��b�he	-������_��N7]�;��8(ȝ��U����*~��[�
�{�[+���� �4,�� ߙl��X���4Ћ��u�?�.�F�3���5����v[��ُ���i:��w��+yd�����;GD����a�2aK�_cF7�nn{M���	X|B��|kN��r�?������o�[��k�Y)�f�Н,�ş����OJ|�H���;��V���������;��W��VRFf�~����VG�5wq�%$�3>���0͞���I.���#L�mR�����7{�m�2{��I]E��=t�'I���1Yx�{�����[�gD���/��f!�٤��'N+*)��_�S�2�1?쩇�ȱ�R����Efi��C����W$P�쟜�_~�ta�׋�'KW��D��/aD
�r��g�4>!�>�L�Y&<]��&⑝��.0�����M��84�%��$�1�X�e�N�E�^�A\0��e�E��
.��z�eG��+��+݆*��s�&IZ���9�w �н��IY��T�QےirHpNW.�mK �$��h�����E��3+��R�(����ߏlIڵ��=��
���OU�t��h��F)��Eˬ��eq$��ҳ�%M�%�+��u]���� %5�(�J�<���?��
9>Fk,��/����g(1�o-x,�଻}]HF��FË�;��GRl���� z.����,��R<B��(���k���an�g(^�/x����抾�m�7^�}�tphcsl2ܿ����"�X&���$�U���^���S��Џ���X�:h1	���L����F�#�?$ �#N=˩sP�>���=���A�Ş!��_�y������>l��:��?{ �@�;��D���������g�)�����o��{K���6�>J�f���7n�#�������S���2L	X68j�}��U6�N�����+����������뒙�0.!�c���YL�x&*jU�z�ӈ�a�x���_,şh��<�2��=��u썏��h��K��2^������M.�NҜ���e�N�l�H�
lzL�B��)�#�����L�/�˛��
��<,,���|_�τ�5��=,�^�Ҩ�N�")�ؿ������;�V;�����ⶱvB�h:p�]a�� ����t;M?W�e�1Ǽ��������oKv^#2�	�9|_7Vk�_X:p�������������I��U�sE�M�����ՖL��:��^B�����G|;����~c�*@ݖ5Mf6���Ów��o��`p�d���P#�VC����r�A¢��m$��,+X��6�=2�b��{ C���4���{s�(��EŚ?�T�>����(4
<@ƋS� �v�UZ9	�U>f�ֈ�^�ȶu�5?��v::x�D�a�r�cu�I׷'�f�9�����̀(��l�H�=���J�u��1��V�xR������s�&��%8�*LE\�M<UvHU���>^�l�a�vr�S������[�4*��O��#k���Ö���b��[��ޱP<j�7�)�l�fE8�E��M�;m�k�$��}_]C��j�z�-�0��/h{��	b�!��k�Rc;D��P��Pieg�."����1����t�ūѼI���:�g��9+�SL_E�ܭ�f����
�x_���L��|(�����$0�s�9�Os���` @����J�rs��M���/֭�)ne�}�����ح�Ӽk.L�����6��UˠR��>�@�D�*�1�55k.J��'�FH3�qD��F��2�3��aRZ����*�Uب7Y��ޖ?#I��T��tڏ2$g�I��"'�e����t��N,� �f���=9���/d<��%^���ڟl�b�C����ְ-�ʫx�Bu1��;�Z^�o�U��r`� 0��G�g]!��q��;�u���*��"�da�J��f�P�a�����0�JPK�I,�ʥ詂4�zT;us�Q�g�-(@��r�����1L�M�����B�p����|��W3��92,�1�m]]�l��FjA7�������#i��yI�6��tHU0I^��cN�Q&��!�gp=�cw�fX���ٯ:�]�8�y���0�>��Xs-��4W ���4�ď!�R8��|��FK�a&d��������V P���!�ƤT:��=��K���ռ�Ze�,�g�Z�j��TU���nWHjX����;�����1�2�Y�V�������k���� ����O4�3@������Ӗ����{2D���h�#��'%d����`��s��o�l�|ֽ>+���q{��[��x#9��=	_V26�ȩ�S���g�(�qF9�K���3R���<h���P.L꛾5��&3��@�ƍj��k�d*%u����g����5P�^Sk�-zH+ �����v�Y@I�8aC��r�o1�I�)��7��,W2(�)�A������sIE�w�v=��]��y?�B�}�m"(�"` HI*�E��I��Y����%y�_&$�<I��H�}`��fH׍�p0S��U�c0��hԼ왩������~���-��	���S&>e0Q6Y8����~�:�E���`wY1�W 7X#�q�"����	土�������#�H�eDC[��J�va����-��O�j�6㖝�dB�J��ע�h�Y�/T�n}�?�Ԕ��+6�.��E�,�8�WV��e�c�[����^g���V�d�fD"i	(��s(G�'e�JȊ�6�TsgL��9\�F�{�9`������8��(��Es��v�?+���!Nu����tn�T[#j���{ h5yЍ��I��T��Q�?% ��̄�� ���g����ǽ�:8J0d�RD���X��Z '���L���*^쵕���L�gLu���aIb:��cԲ�@���D�՟b���j�Ga�-Ҥ�ơ7�Pg'�D��8���ٺr�<Mu74>~�8ܞ�EېE��Y�<+tu����q,�w'�R��49���2�8'f,G#.J!|'�Z{ê��1��WgQ>�Y�$�&1�,
�ĕ� 6�Ֆ��'���ۜ`Q�n�L@*:���-�T8ۅ�^T1ͽ�
a�ό�^����a�>�r!�?|m1�g����ô1�s�A�o-?��_j!���R���������ڭ�l1�*�#�}6��N�}���<�u�N_�&k��d��y��p�=X�/�/��uoE�f��h~���57��� �������f}]���p��1?�Q�j�,
��7�rԾ��s C��hH*0i�f)�CysC��.�ֈ�z�,�AB���1$Wo6t�
���q�]��b��3�U�u�U�X��V�M��x�ʛ�%��v��0(٫��g��Q�TlX�7���u \~�4W�q_��j"���-3,.z,5q�7��O���	���)Ѯ�����A� �7(��6c��;�2yJG��q��f/7w7��I��(XAŋ���wx;�[�Y��o(����z��d�+����>y�o�s,l����JS�>i.-m��e �q�ue�G	߉u���/_��O��#��g�j҃S�n�J\����0���ׂ���;18@k%�c̬�Xd[�?}�0ś%�`�ŽKT�4s��
&�{��%;�j؋��h�Q*��J������(7R[�>3�W�1Z����ޞNp� ���:�ZU{2B+_>�V�em�@��T��:���I͡e�
�H�"���>��';��|�|�7�Y&���U榃�Y���$�Le��)��kw.�oS��-���+����zm�ޔ��?�����l����C�ϣ�6�$�:�c���/�{�(�ʊ�X㡙��=k�i_󃥞$�*�u�[�bi*`�������t��ָQs��`P�u$Z��f�f`$c�-ԏ-]IP��U3�EQl��p`�!siU4P![�wy�T{\W�����#�Pj�!(˩H����j���?g���x8�z7�ow��o�wy#h6w�sd޲���{�N��X���T��)2��V�wu(cg������]:-Z^�G�&�}�O
%Lk.4L�:�n��1��C���D�[�b��#��R�i�t��4I��]j�Ax��֞���:�QP�zAm<��Av���� >���z�@�I�n����6�m���������UN���T����L��%]�rD�	�:�Jv>��y ӽ׬_�P���� �e��a�Ne��~C�M뚸2N0�0�iVϔ*[(�䰝!�z�>䉇��{;�:+`=m�+͝Y1���ۡZ��LNcd��2A;F�*\�M�=����հ��]r7���\���է����,	�.G�E
B�xg�����F"PZ����cEk�y��2	�[{�K�]�6���Hu��.4��f�f�:����k���5�?v�*�� �X燸ϽU�l� cx9�0���*�u9ޮ���,����k��F/v�Wig��
[�x���)��]A�e��0T9:��*c���\�{�a(�|\����p�%�0A	@q*����g~Ѓ�χ�W\�hn=��<�C^ʯ8�szuةT>�t�:�_s��������Y��/��6N��������^������9��z�2+������A4�8KE��4��z��}��>��i#��$�|�s���BN�x��R�8��z=8�%Mv�0�W�����%{�s;�ֈ�z�X�UL�T�[3���*3�Y�rO��񔄤~OAi�%�d���t0����b4�K�용�>ms��B���8��$vZ�7	!	�����X�Z2�dZ^����!\e�4؉���)B�}Mh�f�tikoh�&=�$oiqoϸa�zL;��p��4�����2e��Gw�X�=�ϕ�FI*K�e �#��l]>�J�Q�.����k����,��}[
�f�����NӔjqx�7�����M������h���ơ���u젴�Q�t @�N�[:H� ��Y�Lw��l'&� ��K��5(��ϕ�e��&��z,�˧�,Pd��$�#���nK�P�6T�Ͷܤa�Q	�?��e񼞽��:W�Х����^f:J�lR���ֱ)������p�����(X�ު�	(�C��-X`Y���ǘ�5t�ю�9�jȘ3�?U�T+�u��4!��8�\�}Z���O���BF��;'ߏ����F���gPH}e9�P���cq�U_�؆��e�Z�bh��Ǡ�du�n~��̶�}P:�R��P������q^S��5QE!�j��Sq{��R���3��f������z2��/^�<�=�20#�Z�}�>����Ks�����O�QQ�)%��L}M��S��F��e��s��������HB/�l=}�2�^����)�C������%��Q�JL��/�Ŭ��v%�Dzpxńu$s�g�F���;��sI*�ޓ��w�p��N��>�я��P7���{K�]r�*z��1"��|�(�!����փt'��� ��h�|l�+9���{轂Z����B�!9����r-��:z�iכ�����a��=�##�Ƃ``��u�x�y�b�R�H��$�I����w�X�wAH��� ���+t�}�O��
�?rQ)�a,�z�����7�U�q��6�����m̢&�l$Zg�J/۰���#9�3����f6�\	��^|���X	*����b� C( 
�M�>�HHu�|f^�yq�"������~�N����	@N�r ���
��*����!�I5F���3�Ҵ�B�0�ciEL>`;�.��q{/d�uXH:�u�%2�<��vT�t?W�A��i��\ ķ�<�Ǟ|H��}���`�����	RM5�5��W��y'ۥ�����$$w�Y�f�� �C��#p��n���+�(��#@��x�B`,�qm�N��ŚT\�h��P�o�v��r�����_ݫ$��=ۂ_OD�#��8
�v���Z�I(�W��P���+���ޑL�3�E�5�čՆ��;��C%�OS��h0 ��,�ј�)��Q���]�I�kl���>�| J����S���jY��/��� #)iV��y��7�;鎕�=ޟ�<W�Ʒ���ē!���{�_�H�TRB+���9m��[16���xzl�N��Z7���M�}���"�g�� c��0 {�@����X�R����X��Qj����
;�ot�C<��4?�]c1�B��
(��a�`�)ư���F���oa�[�J�Z�t��M+��$��T��["�L��I� ��D�p�h���AfomXF�U��J���XP3Ǒ�m1�I�3�J4d��u�
@�;�k��+;J*@CmJ+��2$5��qd�X'���,'qhL&b��i9�5���a`���f�3����.n�N��^��H	A��c���^R���L�ȏp�=j.4�>�ք�-�
��|�n���Q���IV*�yv���
�건����Â�ͼ�yw��n�yd�c,����Z־+�r�A��z�4���"k�R�>�?튿f�C�s-�:��0��1av�����]j�I�Q#=9���L������(�jy83D�P���=q�κ�n�a�(^��^yp��V��f	�eI֩[�z�
%��ӬK�� -�T@�I�4f��X&�h9��SD���Z��!H:e�Z�}�c]0��SI��].aĻ|�d�+/��}�皺��:>U��F%mN�\��_g���q4�1��[B�-�y[$�>��y����ƥ��Xf��u����>N���'9��0��֧x�y[|z�Ob����w'jW���Q��w�W � �Т�s}�)DT��\ycU�\�7����R��T�����)b��jλ�_6�@<a%�u�/~<����'�z"����kt��*�W�T1R	��vS�H�LXq�+�=i�?����k�hlF�W.z�r��ӆ�d��a�f�s~t}����A��;I0��0L�T(gZ�ɞB]�v�ɏ�'��uj�ějf<��w{k�=l������>��=e����I�6�ƻv�s`���M�C4�A���V@��s�L��
�����ٺ��u�t����������[�:���͚�Ո��۲�%dPvC2�+�@���*j�:#����>rFN2c���+o�㼘ŐP6�0=`�75�~�lڀ�����Z�L2�?"�����`lOھ�>�`G���J�k!r�	���h"���sW�g,�,�"�♐�����a�A�P�E&H[�,�T�=�IdCj;X��H�+k�K~��#�iAqe���-knʜį'P$"]��p�@�{m{dJߛz���2q�|��9��I��CSݥ�a|�IA��v凩�ZX�)@�)�ȿ
	&�XF0hg;�]Ӥ	Yl}�`�e�?&��:$��4�d+���Z���7o��M2o����3_��������C+g/��Qj���G{��2�B���^A�#�o5+���p �E^�7Q���R��\�٢�	��2.���Р4dјNǛc]m�b�>���O���Q�"E�Ha�(��ʑE8-�ȓ��w��>�h-�%��X��H��=��#�ң����FO�K�p�y����{ή�CL��̢�/f��	$ε!�~� ��Jj7oU�S�ҿ��'/�,56.��4�9z�5�X����a*���!�����#�GR�`$���x��W��r,O�"�CJkD�~�t���MOI��3k�ߘ�`�����m����W�����E3oyyn]�K�b�9+ڽJ�iD���{Vq����ƪ�̭�g�Nu����tb[�k5�I�Ŏ3%�]oW��2̏�7�}p��t�Vg[�KO���dp�X�$2:�w`z<┅���T��c��Xs�Z+V�t�-҇��"�@K�3��R�]�$��J:ʐT��\�D.���U:���;��YSjN�,`�K;i�n��8|�kL��Ő:��+J�Σ�M��c^�ϲ�ȗ^��굶sII�rE���/&�����e���#���3h֮z�1��6��-�b��N��Kc/B��_�[^��ژ���҄fѫ�:hٺ�Mjc#"]�v&̘���"��xK����h�K��5	�=X�m>Ze�e@�
�3b����䐰;e5���YU��2\��]PR�r��ȱ�2j����v�G`����Z/]Վ�)�c_����Oi TU��4��T�j�K��l��iCg�h���E��F�ܯ);�M&�?Pnh�FH6_�2���1Z��u,h���̵����L� G�5>��L<���.`�/7�lR�)�G�=	$�Ք����uR��/~M<���f�S����m��7ٺ]p���Y<7�#����l����7f����`+ X�P�R'��phX��jxSU��Y�;8:r�
PXk���v�־�gu��D��܌"�qWw��v�QH׀7�e�f��&���Q%f��2P��;�K8(;
|�+}�������S��TN��� C�50)Uk�pa��laH�����t���U�쉹����\��L�X���K��\�׼���7˷�#o�R`mȋ���ϴ4��t��5�K�_[����?����}���t7̷U��ײ&+��i��;��=�:iV�x�"�H恓:ʼh������ #e���~�<������KT�u��f�,���_8�=Z�6���������LX񟛞9���S�T���
�qff��ͽ����>j��aY5b�/-u��*�?%n|.Q8��.�yh��Q�F�]�v��c�`�"e�g6B6G2|z-
l�<�Q�%|�^H�����چ?ʃ@��ż�����2���sC�A��]7����.�G�C�z���-y.���Q��k���H��ԃÓ�9���lS�:|[�Z��b�u���N-���'sh��������XM�`��'�n�N3��RX�zSn�>]�\�L� L2��8�?�������k��꿗l^;�Ѷ��|̬�o�8�1�%V�Ұe����pwhj���P�
c!���n\�ºiў��G�=u�n�ţ�uh�g���"N��G���|�P������#!���K��o�׽�~�	�)!�����u�H�i�RH��K����EQQli�]�yNC;����a�:�;��{s�j���r���:0���7#%J�2�t͗qZ�$=%�AO���a�E������N
V��-�<IΝ��qR�r�L=?�������;��P��~�JC��}�ʽ*.iF������e�U��W��]���W�ɋ4�V j߈Lvߎ����|,f��d�x���DU�������O�F��]��P�`�����l��Jx��(��R�#$�1�oN�Rch�pf����6��Q���N�M��;��úv����/���o���.�ҿ��'�˫c������x�\�ӹ�}�E�,�|�#�+�$9*j��wqy{�U��d⍟�|�煛O�6����,\�*N"V�E�}�;ֱ�%ą�"A�ޤI'��.cZ�k�u��Z޴fĦv�Mww@4p�0�$��D��a����z�2��x�ت��L+qGN��/ٻ�ޓ�l�f�K�Y�/d��4r����J�q�jdx��̙� o]��z�Ray�:.���Hy�#�i��>��w�0vzhZ��t�f�!g�n�q�us�4��Ϊ#�������^�3+Sj&]���e��M� B�۵��+��<��C���R��y*N����xk��e0�\�{�[�����-���)O�P+�����/Q���1�9�k��N:���ݶ5����k���	�-[{�=���6�_����R�w�❕;Q��9�n_�  ��KfF~��Vg%W=	�FJq�	!�X�y�բTq���eCDZ���I��Ky�l?�,�0��="X��ʮ�{�_+�[����xO-���)����P��j/Dvw	���>&j\Z���[�/}��� �=�w��#�*7+���^�h�xco%1�����9%y,����廫,4��&P��)�9VxH���{�k�9{����p�K���u&�Ds��Iga��f��<U%A�1)L��7b��s�8/�_c�n^���S�t���9��1T@���\�+�Ύs����ϭ��-�{q����j�7k�)`]p�N�*�l���Y�+���,8:R�͇ ������a��ۯ2r��;r�ۍ'�v�똺x�bj[c�����;{%wK�߼6Ӄ�70�:����5�����i�ox���BZ���p��j͋&6j���ۯ_c�)�]9*��qccK��	usC<
?�(z~sz��խ��.]�Ѽ���t�8ЂU�/�Tfhu8&�]U����ÈFz���	us���w���G��y�S�����&/
\37�^@�_�B߯Cܿ�j�Q�=�"�\]�H�.����}��E-�+A3n1��@�)Y9�����gש��"s��D���C��0�^s�>��s�-^�}��&�y��Rg�~��j~���S�'R��q�����4;����u�j�b�������8�W���֭�d��I�k�R�
a(����+e��S��״�T��b���۲Z��9��F��#��s��NM��#p �iP���­����G��T�ST�'+us�R6-������Ci2��V��N"kW�Ö�g��e�I��e�y+w��r�M��)	"Yw��n]}^b�c�_���@�~��)[�y���	jiQ��6��y��h����x�k�{��ݤX�~%��ӭ��-�����쿯�к`HX�������C
�ў���ư��Q���1��Ge��4 ���'�d���45\�}��7��+f"�o*�oj-�P�c����� @p�/n��8[
pF
ٍ˃X�E�:&��0�8˽���~��15$�,�3�ؒ�`��A���Jy��Jſ;m� M	��Xb9�/�{}��~�9Urn�ق6$���U�y.ur�ؽd�Hr����1��MX�hj�aAa��(׿����k*���jC7t���HH8�਍|O*ŧ?�7X��O���7���g�9�����t�Ԯ=u#٠����F�Ǭ���J_�W?Hһ�&\��R#��6���}M�L��+������x �J��������G<�_�g��?�����]v�X�Sn5Ƕ��l����K"�WȐ����vY�9`=���<��Y-����C���{a8������}�<���;�'�ud�����=�®v�ǎqE�;�S��I�4s�Ԗ��ʽ���+
���@!0hY�B��ݽ0(!�(互^L4���{I'RIwy`�mak1� �9�'ɽ4�j��|A1���|���	�f���GDX����f�{�zO,�2����j�eH�\XPbH֚��}20/�- ��<o��b�����%�%��Qg�mI$\���(�p�I�h%�U�4F��%W���1����]�Z���Tz�����i��'�	FLɄ+����c<�5l/I"{�"�f�e���@@�4g�i�	}��a����盀9w��5O'n�&�;����z�Ԍ�����۲�N��+v5��
���n���N��8:0�d�F)Rb6��;�ڄ�է�������H�y�V��͓,��ws�D�$��AL11)ӳ��x��k�C0g�q�����B��Bx����S�i�b�ț��ԧ%k��@���e{h��֭N���`�-̋�6#ǵ�o�f�d)�a�{U'�ֱ�&��6H{<�w����zlNʑfZ��n߂�'��f�����0���Ja���ܽ[���"��5갶�;�(VRyz���NO��ǜ>���O�^i�VLJ������5R�Ꮮ`����o)���-E������ւ&,2�){����; I��m�Ρ�~_�ӌ��Aln�K��0M�S���ip���H�Eć/�%���M�8�~�k_W�_7��.��5�#����D�Gch>�r2	�83�eB�@�2���;.[� �	��a"�����SX�iұ� ��ܕgک�d��^�٩^i:QWM�56�����!n��FY�Z׭��#�#��A�:�f�)���0��,}=�맢�yϥ$�\�p�������x^~q� 92M~״@�r�S�N���y�Z(�hy9O,������T���چ_7���;5Dd\�uXQ��B��"�n,S�Q��S���?8��.7�L�y:�w��76b6�L ��Ai���yj�u�yM� ݊�t�+�e$�P��z����\��/��"�C�<o���L�L�i�
�����Գ�I�졷�xE񚃁"��L�7�CG"Ƙ�/>j��R��M��� 66�`��&��r��J�〴�j8�&�9.r�ek������5����ޱ�`��PZ�"���K<�� "�Kc��:��K�P��,c0o��wcA�A!;\��ӳ��]�.�.�W�.k��t�z�����'�(-������/����>�9f��ڢ��Z���̟IQB�g�.��gE��#i�.?n*Vi�X��ox%u*Ȅl݄=�Q�*k�lfu�9�r8H8��pUep����,������֝�	)K�>�q�6���J{ң|�GKq�L᭒*E�_c�6��_�k����S����#Y<��AE�*��V"	N��dI�&dge^�8Ԥ*I�|95������h�r��/�O~�r7��`�D;/��$귥��]�AJ����,l5���R������%{��T6�M�j+A�#tsG �GfG5(X2g+�����AG�~Q�����A^Yڡ<Ô��A�>����"�j:G�gc�� }څ��S3�ҝI��xԆ�T�#�P�.�����������AmB����r�!���+��t����ĝ�2��W�&p���-f����JV�=ݞ��w�N>Q��P��������w��p+���ꕗb4�G-�}@�À��r��]b�}2u�f"uj"�[�[W�ˮC�ܹ�U^I�ڮ�殖g5/�������}�"����~�����-�K��� �ņ.������?�-��z?J2��^�)+���K��[9/�b@�e���^�z\�9��&E�B��+��?8xW$W�����H:ռ k���H�])��KR���Z5ƥ����'6s����u4 �����s��-���"��9��ċ_Yfk�v�J����I6�8ų�Tsr��I��S��P�ޖ�8e�8��rT��tҹ���������p�q�6�k�36ȩ�,71{��~۸�%���z��N�@ �ay�-5;�ͼ���G�%E�#>�s�#Pc��d���A�Ĝ�M�/�t�6,3W�#��`��=����Az��ow���r��X;�d���w��LJJ�,e9� o�:K�X @���J�ﾈk����ה�o5�&k�1�	C	�CX1kl�)&��2��h����zIs�t���K��_Dy�rȅ��D~���'�N�ACz�ؒ��h�P,����͔[���ŋf��TC���\3 e.wF������r )�+�G�v��nY}X�0��ɜ�[�ƙ�#��G�8"Ō�ěv�=3�O��EPs����
ky�A�M���t���[��Q�� -��Ws-�������(�n�=�����@V�6�o*��C����Q��z�S`&���v�nPNfKyʮ��nN�ɂ��Ԣpi�v�zŢ��I���sf�G����t�AQ4~�Σ�Ai8��F��Σ�h�����n�.i�Γ��8�{y~���s37���O�����8|U*l�}����r�uZ�bY��1�UE�HJٚ�׎�3 E.W���A��0��֖6��@�_���#�#��oj?�i%��i�"�̣��Ё4x�U��M&.M��,<����j ��n̻l��l��G|�{ٟ�6�S�����E�,��%����������74�?<Rǋ���O晅������]]]��[V�Z:���V���c'&��po��n��m����v�c��e;��������[��[�!��4wkpI�����3��3�-u���SW�"��Ѥě��~���� Swg�\ó��7��0��������3�a6���d���4W�d�⿐�w�/G�{l
rV�켽l�/'^}��}Ylo��+�4���*��V3W�� hv�[��WH�\��?쿅{ȓ�Uk������i��b���7�g��MW��������`.����(�mu�.$L�P�*�@OW���M+�\8��#�#�w�1AL�����5��.�����6{��2����aS}=_TT�v��Qg}M�+����3֦�r�g�4��wÏ�?b�qV[
h�O�`�k�7h4�Ь�p����J�u6K��$�9��̙L\}�nC��T��Z�T��z�����*��/V����E_0v>O�so���4��y�X��*�� 	�=�L�a:"7���P�S�עo�xօ�s��H%��d�=_%m���J������}S��H�	���!^!l\�Ǒ?�Tu�~�����؛q��.�]��Ȫ"M=�;�Y������(�z,&�w�y�WSR��3����h���������*�Z���sm{w�+U'��ǛJ'���S���1k�/U3�b����}��8���7N팛���kҎ<�Ps��C۞��CG�H�X%�<�GB�1i%| ����Fb�ᶍa�c������������v+T�)�x��f�*�s��L22�������������@-��$WND��4s������S�ϻ�n�uS���)��ۏb�����e��=_�w���^�v����'���������X/$֟t+Zv,��(6�^hf�,^��_8�pu-�q.Z�Q<�:p�uޏ�g��M����2���k�S�.��&(��c1ˈ'4���kX�Fr��J�E��,a��JL\�'Jkel�9ʱݔ�^��R�.�S����Nl��)/�'R]' T�:`�X�#݌��9#��Y��w�'���*����*�	�)�I�D�6YBƙ����t�D�J�ķx�z����p����m�p���|j\X�#{�"�H���$���6TA�=��9�Ƶy�gϻ�N����ʽ=	EP�ϛ�tD��tؓO2F+h��"gS�-[Qڼ�!�;�<=���[v��3���]���hw�R#򇹙
��1�1���������7�~�+��\uS(_��6U�^V��������Ŕ4aW������8͡�}=ܒ�~��y4l۳�X�A�][ᒆjA�3��|�K�H7<��{����/Ş�1ez�N�P_��m"�����va��=�N�,�����Q3Hql�x�_���i%{3n<����J�`
�W,h7ߐ��\a�A8����È�H�з4����DPp ��J�>�M�y�o.�ax�6��<.�֭�z���;�����=,N04�l�r���W�t�~�2	�2�cذJ�\p_��@����׵m8Já��F$��m��C�_3M�d����������5�N�FFF�zZ2�SA���?j���MEpǀ?a�g}��6/��+(�bSA�_��Id��w�.5���ܠC|��Y!�V66���_�VS{�i� (=O�=q$#Z�� �D�Ӄw�ɑ��B�tT�8��F���������3�s�7z7�'�;/�e��tcN��Q�拁�a�csW��~?Kq:M�	+��w�-�s~6���A�c-V!�����?�+O,%DD��<��>sմ���r6e�4M�t?��AGd Y�D��7���v���}.�����Ş[ᵻܷ���֮�����;�4���͟��4����߽��V/�vy::M��i��	�OF�?����<@��c���Z�%d��QV��=��[�=�]�`�;w��m�?{�i���i����c#���Y�Cu���[0�H:��J��u���o�G���n=&��\���N�{;��&$����}�*G:�9-���އ��S�>AVի*�F��\���b~n�*��29}3�D+F{	f�8�}_��/���Ui\����y��􁴈)����6�����M�?;�O������"V���L}�t^�����s�c���O�-/FW�S��n�Rk=�29�3���Ӹ�O��^+���J����>�P�����,���������$�V%�!��=�-�%��b�ɒ�D���Ʌ-�L�^a�.�eg� U"�m�qq��uͧ5�]<�@��y2fhݏbL�x�9fQ.��/{�xvDb����@��j^0��<J��s��p����;��/�P����'x�&Eӈe�j�������=�ھs�}rO���y���ڇ��1�q�q��P��)�;cg��?�1���-	��\<{�o��"�v�
w�L̇����C�Z���קY~��,����i�n'^���r��־��E���nv6͖���^*ҊP��2fOU�PG���t}�) ���zm��]�4����k^��j@�贈d��ۙNV�� ��o֤n����������o̲B#^y�0���j|&�7�\�J��o^�a��m�3z�����I��X����v�X�u��7#q/�\M�r3?�	Ξ��f�@N�\̓E������a��KRޑ��y�AJ�l�b��ɋ!���1�@���$�r�`1����D��uւ��&�)t���4E���(���f5c�:����b�B� wn��1/q��`���8���Aw� .�_�KUm�j���T��FU�){���w��lv����+�%g��PN$!�!
=G�#�XOfK�G;`�i+�^3�8,ov۟���2CaϨ}�<d`���3��b9J�ٞ�)��@-��}V
��@�tk���r/��cAP7�4i�<~͑��5�A����8��Ԋ,;'l���t����{@�}ϙ6�(R� ��������҄�t5�]2A�6�����@4�T�v����^�������/���{|�ۄ~0]��'u�`��9W���"��z�C���G�x�j����� .�x�J��bY��r����9׷�$Y���� ���b�/��ծ6��x��G�7v�?����(_6����/���
���G�3.�N*:*��LL��XZ"�j>�c_U�s��P3	�c��J�gF�����Y/ڞ�d��R�#/������Ǌ�*�0������퉁��Ө��l)��S�2.��+q���j�޺`�j�Tk�؉f�8��
��M./�\)\�6�Oم��v��Y���<L�A�rJQ�ն�xm���Hl�̠�3�h͆�Sl��Z�fy�G ��a�����*��~��h�SR�F��ڴW/�,J�T��n�6Ѻu�$X�,2 ��F�R�FZ����M����5���kߜ5�ě���PI�L轳�3c��6G�������ڕ,��H�pޑ��J�P^��%%��W��y
��qI�����8�r���/q~���ʄ9��	��"��4�h��ǆ�CU&d/�0p_1`z�^����rmW���Y��3H}n���N����Y�I��w�*+�;d4��\-]���ś4Z��9&���7����=�seЊ7d�9+DXRNߐr7����t}v!P�2�R�6��dj[���C��0�M�ӗ����ȶ�?�_Y"�[����ɷxMO�i�L�_�aȃ�̡�_&G�g�����dվ���x`\SXZ�ɬ�_^�qu�U偡�vIwOH��o�~��i ^K)�����2|+K.��Rhn #�aՍ�OY����:�?,��^S�'��$�S���:'�T���1a���q���9n�&CS�|g8eq��9�]�\f̎gS�䲉�,��F��\�X��hGY9a�d��i�?�j�lf���7��;A�#Y���s>nͿMQ`�^y�.kS�HۈA�ﴽ�S�{:RUֶ�U]]%�j�y��尣E��Am*�.�['���tu��
��-�@2���GƯ��Q�iA��p�y�
g��E˪�]C�o�Ls����K�.,�h㯽��̌Ϭ~�
�g�E2����"%�}e�e�dy�r�������-,��
��VZ$�5(;�,��i4��,JB���9c����زz�H�F5��>4���	-H��z�&��_	���z�����1c�5O�R�#NX"���{���S69�m��y\ˠK�-�Q��x���\�Wy���(������޹��\��)�g����ڤ��^/�<h�Mīki�`�=�M���Q�8Q��7����*w?5�$���5��}�͑>������ȁ4���p]<%�[�
g����O,� �'����-��l_B���{Thߵ6�VX���?:d��%���囋�H�v[��sT�#'+d_*�
K�R�hIǹ\T�~��ެ�L�e�N�f��Xg��wj6"���)����q��:9��ջoBt��B��GL���Z�b����x�}t�Oy��8�)�@?��{��T�[Ի�jǑt}���B+DoK��Y̜�2�ƭ�������f_���}>�% �ܣ%�(g6<%,,K~�H"n^�B�J�r���;���I��P�L����U�>)�<���]���A&&��i#�-;E�(��n�U��K��7�����V��g�� �F㈰����T��wY���9v� 	:R\tઋ_�<�ǐd丁vDm���_ByJ/o�̏bkc#�̷ͺz�^5;㛒�m�a�Ά��Z���_lJ�8��-�Z���xW����|=�9�\�mDN;�jHx	U�$���@�jU�{n&ɞ� j�`%���L���0���I��q�>��;���"�V�>P�
|�r�(�p�r�����1I�	�LH����_w���3Sj|����c�:j������F�t�� ���&�`�"W���W��	'����!8�B�l�Ŀ��~}v�h�o0�M&x%BTA;g��Q��bBe1l�e���G��Sa�J�aV���dʪ)ĭ]�b�;��"��A/>��|+�j���SJ�c������$��=��u�S�hD�5�Gk��ȪJX��Z���5��`��&���ﾒ�ߩh�c.�Ҋ��Ɔq���`��0��?�_�if��?��EnI�
kِ����-�)VH�m�e4Ut�y���a���� �	<�����d%���Kәњ�$�CCa +_&��kQ����^z��D����H(���2D��].�-�Kx�գ�;"��e����E"t+#���io��8v҇7ʱ��t�?N��ч.v�����^�t+��s�NF����
1&"�Zd�����κ�=^zg���J��y��yGo55�Q�ؑ7���f�%���=sZK��E�xn�|94��;h�9���	8�E��'.��"좘k>o�X���d�Pv3�t���@��z�-�yN��t��V�ڢ/�e�������q�;*��$�mNn6��_�8~:Ls]�����5��*nV�o�}ӱI�{���h\���4����e���t(o X������k74⑩��A�J����S���;�<h�/,�P����(��* ؍Ā%hQ�*�E��'���]���s�`�<��<��!��a�l�K�����)�%�Y��R��v\�	���JѦ7q�Z�;U��Ͻ��a��+JI���'�e.Lx���a���wc��#�.�\�u��8��_���,,?$F�$Yx�ڒ��С�XY'~�@�`)�3�fl��9����/�>f�.���[��J �q{���(\�zU]�1T*V|n��1�j�y�u�o�dx�����J*�C�m��X�H���!�S�r�r&��f$t��L�#H���f�ɵ%i}���rqI�����Jt���{����(۴,m�������k��9^:���[�)h�:���ΚI��눶��q��/�E��`[�{o��$���{i���*q�"������~�aos�L���-.�8��{�\�|X KFB�ǭ�UK`�ɔ����A��|,�3��MW���u��X� to��N���j�J���J�#�(��IÉ�"��e���]��~��㧶h`�#��L(�$)��L���6�O��2���r��h�-�g�ΰ�xY{����r�Cs���%��"�ȰAM�*V/�;4�V����ML,t� ��>�p�],��]���)��<'%�
e��}(��po]����,�B�V�����fL$Mdq�I��Z�ȣq�onٌ�Re1�p�i^�e�l�!����J����1�NΐJQ��о�l�'�d�P$H�	D3�n"~ �W��BG`��`�c
���W~�x�E�ؼ�ii�����x����bʱD-
����WRe�T�Z�K���}rxژ}�� tA���w�)F�x����R�7$��	�kw���n>���05/�7�2�2����j�?S�ad�2)�G��o�򔌽Ӭ����Y���	o���ng1HFO����Z�[C+���Q�Ob���nD7�x�B�%�S�g*�ҺX��V�er߶Q)Lc���_���MhwD��z���7��;N`L��I��-�R�8�{*����nj�\l����
��5���?����.�V�v2'�R\7�ݘJ�Hz0����}e/t��X�a�e�BK�2n���]�w���b�B\�6�O�4rX1I����ܡ[()�i�Q3+e1W��	����e"��m�c��n��G���I�����C�_P�~NFR�(�޽�4�6� .{�$�{x4�ʂV�)J*m�����s&�ו+���Z�����.C[W�����p����?�"�9M��T�M5RD��צ�#��%�̲�3�{��O���������V�v�Y(�JB+v����Uv^L"��&BZ�Ϣ�9��7S����#b�s(�@�ͭ�&V�TN�iN�^���f��zpH=+!���O=T7�j�h��������9�|�B���m��Պ!��CK\��[�_]�2�	����j^ �׿�n�0>O��5F;����`=
kF�jR<u���a�o|<�2 �u�K��zx�f4�܍h8ä�(��e(�qf��k���"�;�����ܨ�Iv�>���oo�����(1�ЉgH�lqj����#��9�`����񸅊4,4����w�����f)-R1��T�%�}�ܬ��Kli�'��Q��"$�Q���nv�E/��������Y�����3�\���D�#���n��݁��(�]Q�~Q\���@�\��I��1a��.S��u�D���7�Q��m��^Uu}��/���t"2�m��e���-��=���\'��D-��@]I�E��o��С��Jrԑ`��
��;���f𷢻�E�aG��x�rI��B[劈�:�� �@��D����#��DL�D��l �;��)��#�J�%�*f����Q�O��ص�QY�Sb���5Gw	}�9,�a�dQKO�*�Ü�҄���)�q\��ķ�J/��O��R���v;=�;-�j��TY]�����b���> �H"������t��G1G+K׸��"�ɪ�T�?li��S��4��4{�rU�u���0ՁS��r�u#"�!����n������4�
��3Yd��"�v��Ofy��I�.$U�~4ƛ�E](��q�ʇ ��͋�TKwD�x���i���=}*b�z�o��VRD��0x�@��~-le�Q�ul��o�rG<%�Ղ�K�x�N�Ժ~Nl�KO-�ngt�7�t*f�	[�`B8�p\/�w�e��D\q��0��[��D�����"�^)����M���܉B����PG-�P���?�$�l����oÏ�r�~��ꏃR��o��A���Si���<@�����{��2V��/c���4�Ldƨ}>i�"�Q&�X�?H̤-łM������,pq�;�"W�
Q7-�#�_א|Ph��f���zFre�#5-0�m�Hu��WI�@��L1�D�u��	�R��=;�z>?w㻌�߹�9>lT+�o���gZٱ��΢�'�@YY@�dZ��ыzfni�8���Rtf=m�jK��C��AR���$g�g�'o->u4�!�1�7(�W�o����[�#��H-��O�P�!+2G��R2ԃ�F�}��?Z	�B<��Q*�kS���|�u��)&�J[�氂j����]\����$c�;ce�?��&SnT��d1aCk�shɱIu�P$ӫ3��ow~���wB��L���|7�����U(���?3+T��p/�h�K���ST���1�/�en����l��ڬ���lɗb�P�Ʈj~?Ø����CY�����̅�t����}����<e=[���񗮙�)g���M&��V�bf�i�l����ᢇ�e1�77_R;�V��`l
G!*`%�.�Z8��6�Z�5�{4��n�.e�{Č�d���֖��c�*q)]/�9���Y��e�~u'���
Ƶ���*�I���q�Z�����^/c�K��� OqZ���e�Z�I��+��u���j�Q��!��%��	�;-�Z�u�
x��!�����
�;�� K����.Fj���=�{��b
��+�؉�Y|�j��m!�0��*��<D�:Aτ糥��>Oǳ��\��ǖ�����;J;��=�SĢI�
���7\�A�B��٤d�2ESr�_�4?��+����8TV��01� �RJ&�1ȝ�L�}*��خe/��b��W.1�B�P>dӋ��"��o��Mѧ{�c�ִ&68�A�	�.��+�ڽtɮ>9v[��E^<�/o�F�~�h�qfU-����`�PYf��N��흑��?����_i&�H���������z�
�Y⴩��JS�L�V|mHrbнʣpGۓ"O�؂�f;4VR�Y~�S�~�?�.m.��{��A�$\��1�q^z����xmDJ
s���[-Κ�>x񗥱�ך��5��uB~�J���6}�t��쩭-YJ���tL���n��gF�mN�5? ���b!��BdQ��'��|��Z�~G��D��a����(#��30D⺈wiC%T㓈� >r�`qBU��29>+cd(
!��=od�K���q[��ɮi�|5|%JV)�yH�7%,�51"��x�25���0�N���s�oMV���~�#� &CF�h����/R��{���]�R�)j��[#d�q���[ ^�qy��a#R�c[�#辒�Z��8�-�G˒�t$�>?���L��D%�\O���5f�)�������UFMKl�)���!�8��xϺ�M��7�.$1��h���09SČ �.��;�ޫ�����YOY�^tBT�~����xFF���0m��}�,(���oo�� �߉�đ2����:G�n����4�����5a�i ��*ͮ��P��F��x�h�c}�3�z০����I,��$,d&@r��v5m���?�>���0)GAP�re
*C��d�Oa�Έ�Cv�6#�.��{Џ�6�l3��a���B�'�1%�A��,��h��	O��ydf��[2']e�Wr[$��h��0ML�ݝi��������S��=_%���_c�q�-;���|q������i�4����o"W�A��B���L�17����م���L�ᐋ�3�Rr P���D�J>ᱏ}�hpA
�q: �#����?`A��VD�����\(t�R�8��b#QU��B3,ӗ��mZ:d�t!�x�H؂4�і2//�e;g��H�Ӫ����.�EO�m����r��T�辘Z�����OB��7�ї�$DpHV�0�B��뢿�h{:2�$r�����o��ZS���T����@B� CI��d~��9N"/�kF�:^���·[6ULd*D��q#�<
D1�V�u��s�f	�0��_�"g�je������)��N��m�7Dm���adz����~��Hc^�L�� �IK	i�S35믒9~�ʺ_A[JT���G*��
�㷸������q��Z'c$������T�`�>�J�b-
q�Cx���j�$&��o/��Ada�� �mw�<�"M�p��!��b��F-&�*{E)�V�g�=G��:��(n�ͽqd�Ds*m�Ov�����F �V�56�KU��#<���&��9>��7s�hʮ�~ 4���9e��NOL�5�eFyY�,�f���
,�V14r�Dv�H��q�e>�j4�ηM�Pt|\���ݾ���Q��@����hh^%>�x2Ǚ��U�M�>j�U�	�>�s�2�a)Ȼ}<��OL6�_����?&K�E� �3�^�:�?;|���N�����ڴ�2g�jy�Z�n�@٣��?[`
��9���H�{���bU�6B����H	6���#�6�����;0���*��'��y�`Ƌ�����6�t���v����	'�J��$S�����k.���B��P��&��qo��y4�,��=�Z]��B�OC�`{�����mŒ�IO_ S���GP.�i3"�ƶ�����wgi��#�W-�g�d_
�1\;��xk�h)j���X��KH���|zU�hj������:�厅�S>�t?B��Y�z�����s�T�O�T�X65���V������u^����uF���Hr�!�0��g��`A�aR�D���!���D����ϧ�H*O��mOd����7G2T��#[k	�d�W�[+tPGP����j�(u�Ν`LS����Ӊ���j���ŸH�HU�3yNU�^%i�"l+B?��7A,)"����k��z��ǔ����	O�*~�)B�z%q���~��H�`½Q����Ś���7IK� Ԣv�}|�=砾��j<��:�8���Xuh��H���ｮ<S]�O����ў�,A�@��?����b��A���T�N�k�e/�[�I�g(�P��JN�⯋U�3\���_hq�8�G3i-aF��"�;�槎YR�Z�bs�ZEP�/������R�#�a�K�� �#VK���1��b8�?d�¦:��>=���ҾZ�`��*a��x�CEPm�	�ֹL��睼o<�+\]��u�JH��eqvK�UF��BZ�~������="��a��@�Y5�����3xK��Yd�zK���`�Yiv&�yC(~�4>"��'i�GqB�&�f�,>n: �V|J���I���y��b�I��A���A��H*�=��O>�J�u�]��.��U�� Pb�*�k��v$_�Y����`�M��h�|E,����J�d��dy�SbX�k�V>�ָp���v����%�Օ����+����7͚o�Kt��(�_�T��g�`�?ǶaEA=��$%��FX�������ŰX��'�SO�V��ti�co&�Ƣ��1j�d��*R�O�����?vMiرG����?�6#	E�ղ�q��tm�	#�P���/!C�lL3rȬ$��g��aq����4P�y��=Ltw��c�޹�j{vaXT��c�/ū�Ҡ�:��S`�����y�������N4S:@��%������~���'@���w�0�zUe�\�0<��=?���E���
*f�&#�qzWg|���$Ԉ�e)��H�\"�āc����G?2I�W	d�#)�%J���u�&�oyP�:ZDr𘾁��)Q���eƏ�#W'�j�?ي�L�4ΙU���%N�V���R2�|�W�O����ђ
`cR�ȿD��n��}+�rBE}����j��)���u����V�k�F�b�(����U�W�+]�Xp����.2�C{���4hsT�[+h���.����x<�_�?
���b��?/��,��5V��ܲo^=h��|�D\�#��6 i#�o�C[׮�̟��~N0"i���{���FH ��m���y 1���qi;
���qx*J�#����,��x�0�d�a�f�;G�|����.�u�xĲ�'WNZ��J���L�Cn��iu�j�s�+n��%�~�G{�o-��K?�n��fk�'B�q����-�qd�L|R#���r��%=o���ʕh�.����)Y̨2�<x�_o1j��cuA]B�J��nJf������_Uh��HR�`XX�嗀91�$�b�����h�.��۹Ʉ��Pr��u���򑻩�O�R@�K߱��ҟ�����]T�{������	��'��H��g�X�g¬���q@��N��>Ν�t#[j�s�
��w᧡|U�>S���@<q�3����'� ��&7��R����o9T�A)�A�DB�s>��w��ڥ'SS����q=!�}��k?#	u���^;���$�g6�Y�xl�jܸ�hHً�M�~ӷ�Jmc��Z��d\_h6�{����H�����В{^\�ߍ�ŌCs�����d2s�'G��=s�9����I�F䑆��{B�I�j�q��O��}��SQy���Š�c3��ٜ�ڭ�f��~	��7#��XtH�z�X��PV:�-ݡߛul��q���-Y$�k�MIȖ�Q�EDx���p�`��7̭dI{K�'��V����x��>���%��c��Gkd�y�a�K�<�U�#�����j�]g�����a�������HZ���6�m_�3s��3g��~́�9nj'��D�񱁊���l����Y��7{�,���Ş�������|�D�x��{�'���c������Җ~�PR�4U�]�h�;!�_!'���7ua%�L�~�_����)���m�B�=��!�ӄU��Y�zOܸ��W"��y�o�LN���!�==F�;���H`�D��~��T#h��~�9\���5ͼSQ���(�������Z�K֯��KK��B������p1�=�={�H&�kRbƷ��*�!DE������%i���Rٖ��+3e�T��9�E������j�Ƌcp�n���|��p܎���@�
ސ���ޮX\����1�����_Ge�I҆&ASUx0��y`X�~D(���F܉�!�%� "�ׯ��"B�!��e�ZX���Z�����8��?.�=�@�k]��#�8P��s�Q�fo\�"�Ca��=��S���w�������SaMt~����e�Y���$k�$�Ϡ��W}}$����W<]KM�[ɣ�{���ï���iS������E��(DC~R���L����Ƴ��Ʈ���|x��+QH�����"�	r���dپ���*饐�|��~?C��{F=�����q���i����~�
��� �v�?�D�~��c��}�	�>�ǜ>�Om��%�����*�)��*Ħ�f���9����D�hY-���\���dކ}y�J�A�ʰ
���-�?���P�@5�9!*����Q��������L�,�e$��^�B��'�ǫD��aף�HP<�KX2�c��ˉ�?o�=���ey(E~�Hz�A�\Ŀ�*�ZJ��hDN���u[2�8o%��N�f
�uTT�{2���c�]��~`�jQ��{�b�O��YM{��%|u����>���F(#��ِ�u�����%�����r"tpʎ^�P�c�vXt�#�Xx��U�40�Xm��7����y1�+�O����%�� d�n�Z>�x>�j�5R�r�Yu��,[P���*�g�!9]�P�]�W�ԯ�9�n�f<��y��(��hM>U��v���̼sfI��8��U\���2S����R�9�d��7\�7��	U�qhb�v��ϋ=W����O	��Mp=�(Rob���s��͐��k�����
WI�{.��aVz�f_�,.&i�Ԝ��Z����Y���b�w�^�	�JqԷ`vR'�����~뻂���)��/��*K����6bII}�Om[^L|R�7�V*ިzI 9+����� �_��9ݩ���U�!�21�]��U`x�����^�J�2_�N���I,��'�ܙ���G&Uf�Zkb����Ψ�zڎe6$��ƻ�x�n>��1��xT�ʸ0��(;Pˮ�$�-;���.�Z�1�@��ڬz�q�Ӿ]f"}S�Z�e�C"�dd�q���i|�5q#�*Hi��Kj-7��Va!��l����ƭk��&3�Z��)ts��g��L����R����Z�ǕA��-j
�3�e�c�A�*�䶿JGe3��h��X,��[@C&y�[s�*MU�H&�
���_��*+(�Ӷy��!��3\b����0^�z.��J!�=�m�~.�y��s���8���8�W�x�ҏ�^&pp����$�#�e�����+p�U�t��w�>��QH��P�Q�K������,���7Q_���]�v��t�����0H/?�m��f���JarE��?v?>Lu]t!N}݈zixM8���z�xі��8���x�c#<`��H�� ��0��x���jG����e'�N�|+[����2�X�B�N��W�Z����H�71�����iD
�J���G��cx~N6�e�����I�A
�u�c�ښz����Oq�Ӧk6H!�0.L_�L���GXϟ$d���Z��C9�;��H�G���.Xs��`�LY�JO��1l�E#uJ�|�|�2����"�e�ܳ��a�<.���0�0!�ͪ�±��f ����F67�&$�'�3��j)m� OGt)�3	���)ȓ^>L�Ii��}k�r����7��Q6Y�rɓ%r��9�ٳV[]��$�"�;®ś�9��j�Ost=%�|��@��f�[H?y�Z�
�������"�JTXLkV+�n�.rp?�����GB�S�9q���=���h,v���y��C�Mgy�%�[Cn^�?�K�$�"ʑ�0��1���	d䞷d6�v��{u|6bɖQ����_��7��2Ȝ뾙�C_Q�xl���@ڠ����r���`��HJ6L��#��u��?hq"���Y{_����<ܶ��E�<����zk�~�"��������NK3%�Г�<WXZY����7A��$��m�敤T�^�"1��<~"O�.�n�X=C�������"��k�|�Z��hQEj�8%�c�N=�Gt`[�����C��fSGz�v��X�i�`آ�d���.��¦��j��k*x.]� ���#� �4�A�>X�U�De⌹�ۮ!dϿ!J�K;s��a� ���$q�P�h_�3fM�Kj1�	�?�i;�<h;�)�3�Y=����?�ȅ�Z�?��5�^>*��oj�-��PK   ���X	�\  \  /   images/898ac7d1-13d0-4a1b-8b5c-ab7066f4327a.png�W�W��%����K`鮥;%����n��I�EV� !݋�t�>��;�̝{��qft�U𰩱  ���"��:��&�ߔ���'X^���  ���q1��w��S2���t���y�s�p��z����T�|M ��)���YfO�����~qv��ّ��v�C�m��� 91��3�,.���3��2м�P%sVOV����$�\09�U,��Ka�����fv�6{{l����c}uu�ڻ����\"�4����h�v�Y�!^����!7�)�Nʑ��[��������y�B�{rrr/[��q�$�|g�Q\P\�_��m����?���Z�|�}�X__�-��pM���������O{uNF����0M8�W-�Դ��۱�茀��4�7�/c���'ˎ�{ƀ������ka��r-�v����}|/}||4�y}>~�w�R1)d�-�uYvW��������kkkW�O��V.nn�� ��|'��I����K$A~���:���0/�j�ڍ>�^�,��ۛ���x��krΖ[�2��������I����}b�t�#���3jL�Tp�f���%�M��&g>���h����Ŝ#)}V�c}pr`�A�W�rm('���� � ���0���7, ZB��{����p_�u~�>55��ŗ�L7u��aMH����euU�򢻋�@q19n�ViFq�{$'��Q2��SGv�< ���Z3?d(9_�S���'���Jߧ�kc���h���dNF��1�;U{�K�����B�~�o��JL��S�d���b��*��+f`uy��[!s^���w����%]�sCã�~�����������x� �r�fr+�T�^����>uMֵ�컁1t���!��Y*��%p�fWD�����Auu�]��E�R999�e���R���M뭡��'�i�=N�#U�LԾ��<�ۯ���g~��d,x�>�-�&Inv]_���]����*V �|�������B��.{��,s5��D���#��Y�]��f�h,�2�@������?@=Y-���犸��{ǦvFϵ{�����eI��<�T�ۮ�?�=����#D@c]�!��Wg�>6���g�T��Tnƻ;� x��ú�(���F�����.Y����֞N�;=��U�v#�Q�EA��� ���o����T�����<�]Ц���P�U�X殎1��ٽ���ş��z��ɿ�eN�]�jGs���\{{�0W�5(���f��,4��S*��A� sIh��Nw2�J�l�ਜ਼��X�2h��3x��%Ǩ�j�L����	!Y�@�G�s��*�l���#�ie�	IM�f�� �����W��D�����<;a�+~"�
z��;B�t�U�ť�&֗ff�1ɭ�}q��2JZ����vj�6q�^ c�Ì�M���(�0E�⇥�<���-��~ �*�塈(-�?���Ć��$??���q�yr!Y��:�	�7�M��m��;e |F]Z0�u��Ӿj\pW()I�+)�F�8epr/a'?�޳����]_А��Y�5�����ff��Eig������G��i�	��7?���y���yVq�]�x����
��1�fs�(�/�s��l�R:-���^(��6?�s���N?���eu�-�&�i�czkH��Q]��"uj�Fz�0��a��5�f�H�EK���c/I{k`��pG��ߥ=n��[����ڥ.w�p�a�a*h4�Vb%F�J�觍��vgc����<n�����a��eG����U���A�5��֊	w)��~��+����i�f��uaΚ�¯��k����[ ��陙�.`ra�AlqC�h����6�S��'i���nSo�'�$���ٹ����WKF~�!��%�0d\��Em�O]䃍��+��qLi�\���k>
;|P��&�Q6P40L:G����J7>0�e+��f�Ԡ���,��{*�$��Q��$h��#��~�i��*	:�R=�0O�!�������d�!8�۠( 4����U��-�l*�L�� ����\���ch�*���bh�J؆*�m K�1��JM;���s��¢k=�{�5���l^6�&cW4|Y}}wl��j�i{�y������Q�S
�	�Jk����rl(@�%ݴ'm�ڕm~�����=�tLV��%0#)��{C��@Z3��h`��[�0$/x�t ��g�?�H�!�B�tV�+61��BG�nna�R���o�^2�J����+�Oic6|������$��,�8`��~K��	K������儃��{(������v�>�)�����'�ςE�\���udJ�HG����5�ؑ\J�M���M����D[���#y���� طt.����Z������C�+[�H�����nK!IG~\���@�#.f[��=�-�#�=	�k�T����B-�m�7��p�������'��9BL�[Xvل��Ԥ0��L�;,K��Rd�n��5���,�J2^�A�+*RR�����g���U�)��ݗU4�����s�c������Fۦ`e�m6vX�t����V��X7��������F�M���1��7?tK�z+~>�\�鑵z���.���il0Ͷ��z�����o�j���W�)���d6p�n��X�����5D���'�((���W�_��r�wu�5��b��ߏ�7{4����۔iA2�x	O��o�ͩr�Alȅ��o��)�?�P���/J��(��)>�-��qQ֒7�������q��a$��7�N#&msܪ��/pѱ3���H굪F�H%n�58��G̮��*�'B�87�����%n�p!=ExC���'�'�F�+�,�2���(w�Q���Y�� Y�XO�Y;�2�����dI/#|�%��z�0%%��=J������8��]�@y�? gnd�ns��O���kI�dv�E���E�/%����@���q�L}@N?:D���,lJ�#˩��fh7zC���[��K�1Æ�5��Y��5�UEd��{V �8�f͙��:P�h9_���%\�}����7�E�P�E���E��1D;I�8}��rO�C��\�&�Z������8{3ͭ�M&ވ
 p�����4�BtuP'^
��/�Q���[�$���%��U7��Ĕ����v�����Z���*�\�W�U���gj���=}���D�hR#��E0��fi�ۑ��>5eY���3viܵ�e�����hA�v\z��7���r؇�ҭM�iPP6ֳ}��=����u����!x/�E�`�%��c�<���,G��
7Ŵl3���}S�A�:1��	�p�����_�ð5=߉|Xj�W-G4�Ҧ4�����[�8���UP@����m}M*�Q�CQ�{�nK+hb�M��զ�Z{m���JM�W���1���7����h��PO��)�y�~�6�{�$U��F 3��U_���h �=�������l_G�R*�MF)'<���H�~V��BI��vp�66.�+up�nf�p�y��ˬ�������%��#Ҿ��� *b?0r�p )�ʮ_FCg�^�u�NkRa�lI5�x@�	Ub?)�Y�����𷌌z�|�<04�'�m�r%h?�c�;�_O��Q��I�F��bW��9`&aL�8�S�I)�P��M�~3���Kx����ދ���2���qc��)v���4Z�p�o��I��	�jk���4��V����V6��2@:\WD�5F%�D��o��پM��g�\�!��@�����[�Qxa��F]����/���mA�zl tG[r,?ɳ��h|f�C�f�xgW���tg���	Q�!� ����<�2���
��S�����uʫ�H�1c ��$7ے�]9iJ%��K��x|H��?�u�R��䥏�~�ꄍ������p..�Y�ܬ�ܨpS{�!N����� ^g5K��;U�|0�.~\�p��Y-8/�ة�{^|�1��жٟ�Z:k�2rc���yrS���\�M�A�ǭu��w{ۗ�)���濆���w��Xw�/��}��6�'�Z
��b�!�|��լ8#��;�o7���i��I[�P}����Ę�-���;ɵ��,�E.r���aUț��j���}9$���LZ��N�����Sw�웩N^7+Q�ZrDoo�n&���.G1`��8C�
�v�Rl~Yk���J?:>F JM=߹5���%��'ב�pB�U����V��Q���&3��]M}��L�؁����Ц@q%���v���ߵ�y$Ϥ w� ��?��unin��}�[C�y���a	t³�{�}�^���T�U74L-��9�U#��!`ƕ4:� fPpF����v�N��z$9�;q9���cO����{�m?Z۬.j���Fw�*�6��k ��A�R  ��N�2Ͱmz�����B�?7&&��g�Q7��p�%Q�p��*��۹M�[.ԉ�xKK�s�4����e��".�1* �0A�Yc2�PH(i6D�w�`bQ eZ�:�tb�y9%<�	, �b�����C��+�a���&ղ����;[K�������`����E	�sy֝�w��E��W���������̃VެGG�S��tך��X�����،�����)�U�<��x���~�ݹ�l��{Sj�w�)�ƺ�a���k������y`eQ΁r^��;J��r�2m�慗B�OQ9%$�&Yj���C��̪0�[�E�^l�k��Y���/'�O@mILdw��h�7�܉2���c��_q�������1c����~��#nY�JB��g&jfE�rP+�" bzC�Øp��x]�U��� �I�����gN�@X�5`/9�䊌,�&��>�<p��s�ǆ���zu�k@���9N�v�o��=�	��y�Z�k�.�>Q���+	�R��igF�̚��T�Ǟ	����<D��7w���vUk��ٔ����*�'��'L�.��-�� q[PV���eOǻ�W�q˒0P������sۢ�V�SY�n"�T�N4@�y�M�ܟi��{f�=E�}|��_��#��2����W/4oT���=B�`H�֙�ɚ��JS:Ed�!e�%`��n���q�v\.��p�p��]�l�(��"�J\𘵾V�v�m��g�B5>�w�'�%� ^p
q�nބx��+��>�f������k�Wj��|��j���o��_�ʈ{K`"��vZ�,�[����=*w��Y�R������i���
��[˵��ж����,�"8�s/�(a���M��;�?Zr7(l��U� � 5<��N5�?�Zxn���~Rx�$}I,�OYQ(���8�-�z^��-$�W������0cg���Z�	ȋ�)��R�dA=͸���z������Y�\�+zl���y��8Ϻ�q�=�����6:8m�R��N���`-�J|�����,��!V#>N��Oq�g_�"t�uU���hX7o�m�i�Rr,L��z�->�#8ÀU�#�	6�s���Q69��&��w~�4�~���VC���� "�����y\U��j(�S�����Σ�Z�X�k�O	�!�$�~Q��X5�fѐ���,�4�#u]�1N�.8F=�Пux���|���(��:'�/C��[<�AVĐ!�j����˧��1���:�
�]�}1��L9�?eۼ2K����l�vr:��{��_�3I�p��P���fۼ	O����(a����w��r������̒I|=�����|K���'wJ1OU�#�AT?�^
q.b���\�kr���͸洘�%�Ct3˨��A�|ؕ��`�� �~�Τ$�-�'[
iXS���J;c�wso�H�=�
�w�HKP�~�^:=�!���B��3'�z��G����Oʑ=<!?]`;
�6�������H�&��5U��,/���P�}��մڢ
3V���\[@�e	O��i̝�KBm]�V9�}22�)�u1z��I���B66)X&�ր��1n ���Ph�ĉ��ۘ���BG�AAa��S}}ɯ�*��I��z���C�;i�F�DV�O�	�GV6F�2<��v�����'�/qK�E(�Wኬ��b>��Jbd<���T<�VJJJis]]p�R���SM����3�rW�����BF���7��!�����x����!w@=l̺�㮌c��*3��ڂ�L�/��"U`�*_�!��?��^�S?�z���I�^E��[�ןb��R�G#��ݎ�]���z@�������]ϣ[Cگ,��j=���j����4ݗ=��ڱ��Tu�:$sy�ab���0d��1�L ����G����5�>9�iزiK�VFQ�f���u��?FSS���X^s��Ja:���?QY�����]ǁ�%��[����n�t���>cd�n���5��e�#n�{~co׼�X�LJ���%��2���W�`�ee*���K0Ȭ��RX}	y�q��/����(���L.,~�{�r�*�Ţh�H@n=w�-�˄M�8�sũ
�Z�1����sqw��5?�mVYuz>��7P\�?5�*l���R���"�<=�j�"���3��ՙ����-$ ����I�7n���b���1g$���i�����9���L/��q�#������&�FFJz3�U(SR�S��y�.��@*�'Q1���X]�./��f*�����'��$::��Q}kY�u!>K��~�K��z6x��0晀k�˻:ݴ�+#x+A�`w7�s�dm��q/ɵ����\�ig �ִZ�$���H)���Hd�g��u��#�.����[S"��u:�
8��k5Б�~�(4�}��iM#�����32y5r�`K���\c���׍���g,�d���qJ(�HDKR�Wuk�WY�
�ym�fg�ؒǽ2SI)W����qȮԒ����+�ϡ�36ZB�!B��V�	�(�dϓ�S�,�g�����g�Ih�Hx��Ȟ��|�b��.8x������+\b��O�	������_�K9f�Ð��n��T-�w�s�Ǻ�奯O�F�e3^�����"X���/)7�z
l�50v^���f� �T��剡��O�Z�'�jJڊM�6Q�PK   C��X o
7  �%  /   images/8bec88c5-4482-4569-926a-ae76def9d576.png�xwP�ۻ�$�H��*iR#�TE��D)�{�l����A������$1l�"D@@�H� ��w~sνs���;��=3;3���g}��z����}�2�m�y�Ÿ ൴0� `( ��8�����=_XW��K8 �_������" �[�]�S�1����B�{�o}B�/�ϥMT�~�<Ϸ�s2+��&���Jx���]�2M�m��>�y5�׎���|�&��C�]YBZ���ڸ�v��7�A�����y�In�bn��.	��_��K'�$Rk�5`F&) � Z���f+��l-�4տqO�Ψ���Ke�]��g�s ��5N/O�P�W�7�OU;�����W�s-�Fk��"%����
�� Fl�@9�����7Lo�xdY�!�b�'��_Ò���Ԙ�	@1D|����CU=��Q�>���û�kE�f��Aͮ��9� pk��ց
����f�H0"?��$�����9�&^&T���X+NX7�+$��������I���3�%���Ї]3m! ��b�x;�.�@���fa|�Ͷ��!���CjM��p����)mg��{��	��'|�vN�Ȱs�1�B��E� =�աAB��Fh�y�
�i䚶wf�/��G��W��'��<�h�"�b��C�T X�L�M�B_ê�ㅶ�l9?#��:�1��-�Xs�v"�ψ�����	V�w�Pip�)a֌�&�<#r�&A�H�.���韽]W?'"�wNPz�͊H�<&�m�z�X�*0V�s���� �Bw�8@J��@ℏ#5���N>�)8<�|@��m7�@�.l����n��� @`g����
�
e��_�^�� +�����")��P n��P���������
����o�%�&�Cw#�_�?e}ʷ<���x�ȍUPE( @�Y��&��K6�wQ�7��J�3TdQ�jt���̨�9+�ھ�K�*' ��>l�����a��H@��@O��T�M!0��������VM�|8�.�)\ Fu���꾺�Ȳ^�7���wT�"kB���=��P��7�yp�"db��ݧ�Ǳ#����
��=�"��,!�$��ui���1Д%g;��6UgT�hʖ�+~���+&Z��|�����, ��B$�`�"Y�"���Zi��#��ۅǁG->;�<�21@m���R/�X3s�P��鳫��(��T=O���[���ק��A�x.��|G��T�	u
u��x�I{,�t�'����io�uq�-�!��s�:��⣶^��^��G��#��<�ā��t?��z��*�������e�y����=�!9��o2��q�(}�������ӧ{m[��]�M��b ��~?�it!-(�o�]�_@n�|>	����#�i��1<�$?�>Wx_5#�GEV�ϩ�Xl����߄�������B�P�m	NI���Y��ߣҠ�nVI�g9u����th\Ⴢ����c��C� #�y�`��,�m<���Ě���k����z�� 5��-d_tV_��_�_ia�.��42;�wxx����J�*�o�q�:�g�ڶ��TN�L@����l84��"�V$�iU�&5 �'����u��B,8+@C$�+_���DP���qWY��拃��Ć�\~���0�c�΂��R���x���%�w��)#�r���]�lbM�煬�@P�ո��yN^��M �kDpUs�
��&x��0V{�B���g�,��h')�rV�׸���R�ٶp ��ُ���N���MN`��tь��Aft�����"�>$6�fs
����Lp��� ���Y�m8�[�N9gs!�"��1�!�c �ZO�.̶�:�;'��<_?PؙL����X@sq0��$��5&1��A���]U����P(�ܼ]�Fק}[�+��g�X��PBÕ�圬��Fg�����n�`R
J/xC㏙�cI��׫h��£���5ZñB4@����wq�(��M���*��GZ=>��q:]Ye( �l����d�V��R˽���2��u�{
�	���뾸%w������h��|0�3�ɉ�/�J�i����>s��cJc����P�Ye�8ʋ�3*hP���l@.r��]f�Iכ�'����S	������E���}۩gz�c���W1��t3��n{��q��待��K�AUa��U�������쐊\�������S�U
=g9�����c9z&��PY����yiXs�\q/����{jѬ��K,��g�����36�A*lե��]���|e+�^�ǍYf��y��_���7w!l>��^��3�Mk�]2x��(@tѫ�k[�D`�8Q��&ͫ��_/x�%�R@��`s�rg
@_׀�ض���O����N�Qp�d�+��)'��_�f��'�+Ƕ�0+tp�2�	x��Sj�?)/J�tFm�h�=C~�f�����7����O�ԣC3a{�
G�o;���3�H��K?�TP�4�NM*WD7ً9\pj�Q��8i� ��Q~�LF�O�W����s���8ɓ�Ɨؕ��=�%��?s�N2*3d��#R�w��L�.D-���n�މj��3�e�ye^�Q�� %��#_ZgD��z��ٯ`�!x��e�t�>$��BR�4�& � ve�&\x�m�
�4h��7�@('�s�"�������vh��{k�*���>��Ц��q��I����t.D��23�sj�v%;8p#>���\�G���)��^�����*�-�\���x�7����=Y�2GL�Q��V�1�
�c�����e�m=AK�?nQU��T�x�@�}*|aiwWĩRBJ$v-`hS�<��oz�Yݎ��=%���I�kt44��#Yh�Կ��n椓0|�|��Y_���!��Cg��.D�pqkk�O����]0�(��S��<�
���>(7C�FK��1�܎������/.�F�*s�"IA�׉�6�*����	}��<���+D����¢��'_إw����X^N͒6;��q�[ך�Q�U�_�+�t4mv�:ȋ°������{+	%� �{��;�oB����l�[�j�A�|u���`���y��y��g�98����h2�;y��5��O)���X��xi����Ԝ�o�?M0�ń���UUU-�e���
�lמ��D��=�
y70�Tu��uA�KX.�����'�w�+��݅�gӳѕ1�7W��M�'�vrr◃��1���eh8���rg�Q���9�P������3p�P͇���[}m��Z�,G^t#��s�46zK�R��KQy~�-����`)��]z��6z�h|�ƍ���/�>:�%�s�����f47S�G����k�ݛ��+��88/;��ӿ.�SNx���
�d�y����E�BZ?u���� ���f���S�����#
�z�8���R/�s��T��(�3��\��%.�w�?�f��>upjY^�~��;��R�3�I_�y��{W<�,�E˨�KYq���P�SkkN����Ƨ��,��-w���IԢ��|wX's�TDE��'�I.�r���<��u�������e����%$��'l+��.ɫ � DZ]ys������Z��8R�P�]�4��A<���82���ؾ�av��
����g��1e��!����Gu�β<p�@s�vIY�Kk�z��F�~�ǏW�	������&��r��=��Y���_%���F}��a�p�$g��^c�W3;v��+����z�'�Nm���<6V��b�&�f9}��͊��7�PdN�g�?-�轛�`YT���Ᏹ�7w�X,��R$cV[�o<07ްaY��Ow��8�tҿ�c\JK
8� T�&�'ed���j���3Ť��:���{T��!F�B�dK�T��'~�6p)��V�$�k��Ļ\v�2�0R~�������\�,u�f���+�]��K�.k�/qX�`��4{��l�G�Gpr
�y߉�|��+���E�٦zsנ8��0֠���2�O4�}���؀���Tm�����������zo�Y7\�æ~/���bS\���BvEZ��:�<������c¦gK��i��<[����2�	`��v�2;
a�~?��}bl�$�R��'������hU�b=Ⱦ�YF�Er���Poa�>���?�BŐ|��֚��?��]��,�	B�Ox��&$�ͼ晧b�o~�5�h*;��Gr�-S���6x�!� ��
��p{�#Ѣ�U�@:�#rt��Q�,�|��6�N��\V�VC���
e�d!Q�iT�9�h)t����C_x���5��_ɚ�"^��)�8S�������2W���Cj85�Q����K¹��[���{�B�7K:WP"H̡��৏�r�n>��:�H�^RoL:'�q'�8X51"@:�@{hPZcM�){�S0R}uy���4�V��`R��C�ӑ7�\��e���־�k����(IzC{��A�f���C)m��o;��o_p�jl�&�v�w�Nt���%��c{���D���(����-vv���5?V�9[݉��f��`߭���g��pԌ�e�&+���A:/z +�?ku��q�ۃ��r�u�#�ZG+����tn����)ق��V�T���m�D� �����@���,�f��S��F��Mdf�Ih�9]]J���c	��Ws�Wbå���e$�+LVL�i�L7�()�i��e'z�z^z۠)	-D3����pq8�.R>|Z3��֙����6�a5�"e���2_=��@OS��"���I#��W4�¹U9��2����H�]�x3�$�yl���LΘ�
��U۟�����ɵ�
���q��WZ@�Y��pFM�c����ux��)�X�mx2�ȯ .��]��[�;�H����EUS�'��z4�RS��m�Y(��<\8�"*�$)����8�yq3kT��~ޏM�Bϒ~�m���2�T8I[���?�k�/��l]�T�q�ߟ�|n��B}�ge6?��	6�Ԙr�������XJ��<�f7��\�q� %8��4D�ީ�,k��fpc���(��zFmt��[��&ֵa�����>(/{��]�����`���B���ӣ���F�w��.8��[��Q���,;C��z?HF��~wJ�V��<��;��D�fZ��gë0�]y�������y�-N���͓~��(-���`P ���a-�vlR�w�?��Z�H����K�:>����V"�6T§5>�fJ�m�!��2�hܿV�!М.K!f�D�<�H�!��{�e" <P����t��Ƿ�Jr�%V@��D�tN����9v����A�	^�2lt�D��[ Tru�O�[�Ћ�a��Ӿ�ǔ���ޱ��qtG�,)��qU����D��G���Ay��t<u$�%OUg����L�O�iI%(��	�7P���X���V��я����k���v.$J���еo_��Fz��Fs�e��m��<�}�ý�ڲq�!v�E�E�k���ú�}�ĸ@���Q]�n����/���Q�[�|];zPi�J���g�Y�x���':zRq*�w���_��z\�2�n�c��3>���g�#%�g�t���	��[��z��2 [#�bݯ3�c��>*g�9�I���[�0��@��d�[i�>:-?dv�^|1��~�#H}烪�����o�ԅ��w𭱻}�����]��(�6ÅxJ1˵�&���/�w���'k8��;y{�q#c#�I/��D&o���n�%��gs�~�7D)�]�x��`R���/���q�y��1�C<��#�p���4%)09�҂��a&����|��NX���U� �h��+�v�QT���U֖j�_&�V�������e�)��c�v�t�K�wx#��B����VH���I��j������Jx�m�J���)��p)�\�E���|� ��b,���d6
�޲��"����kӷ.���:CC���%�!6�B���� ;_i�d�~���?�9<l�v~{rAQ��#X����2�H��P�{3���}Xr�d�����<��E4Ƨsm�l�18��_�>��<7֖�,�>n�B�~���Q���z���e���c=�Fؑ���S���|������L����2a����D!@f��Q�v���ؙK��;���ۓ��@j.y�����ۧ����TÕj�T!��%JSJ���B� �f��*ߍ���J�{mկP�Ql���>'X/�P�G8�V�~�BE�=�c��턧�r�n__XX�S(�8h�a4\K���f.���o���da��K'O.�0�^c�Z-���t���~��r�����BfCx²������M����Ũ�>
�G�zt5"���7"��h���6��;7�z|��&��;Fc�Ғ����dI/L���&-v%�Fv�Baؕ�fY���)g�ᚸ�1]�|��9[�������&F	��
u.���>`��1�/��0wț]� ��E���c,w5L����`�sSA��;�{N{�>���d��6��q���Yc�;3]=�i�"�rcu��oy��>�~�Q��<l��������r���U�7�����Ѹ�����b�өAdǼ�����V���?#X\���|a�(��+b-����p�o���>	�>9<�>h`�UL~y��*ۛ7�=!B9
n7��kت>���(B}}�S*�}]|�Ɗ��#;�+j�p�*8�I��:�8��Ք/�,�{��vG''_�M�71�T�1�X�˫��bE�]YF�g��&��Wj/q�IF�-1Z"5-T�~z�
��xU�}��<�Xi:�>M�˴[��1��������Y��w�� PK   ���X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   C��X����?  [G  /   images/b3b368a6-ed54-49be-b991-e8c4c6667997.png�w\�]�/����B�&   54�(��- ����R)�A��N�	(J��JH� !�@Ȇ��v������߽w���>O��9s�̙�Μ��D_���f-�G���'��;K�΄ɡ]�?״�c`�;~��BڹG��������������:1��yy�9<{�$��뒵����p�A��}���ՙ�l���e�nc�S�Q��N��~Z�M�,N����>,��ہ7�n��Iӛd��b�>�[��ዎ�տ{/��3���J���s��]8:=w����]�02Q�+�Ȅ*�(�(㼣��2s��A6@xF\���o�~	��i������j'/��8���pR�N9���x|�q��~������������|�_���og�Q�_X�e����ր��<s�A����S:[Q����b��O��
X��T�6�+���E,0�!���{�j$�J���,'��p gUM�Q��5���fTR�1Lf[C"S��1	��ӌ�;?+��G�����
)�e����y�S2ۡBp�/��di-ep�y�<8=���ʩ?�k�|�����
Jӗ�V6O8O��㧀�!�&��!Ì�!�xly2�"�g��ʿ�B��~��U�����-)�4�p�A��8 ���f�kԅ����,�����}5[$氡���x �eRl��D2��Œc���s�u�2�Ox��M��Dj�4��;�ۈ�F�$���]cl6Uǐ��ŵ�L��_�푇���Nѡ�P�w|s�	��bC��Os��s2���y|�����X���z�|�)��~��۔�+� �
�q�q��dv�ݽ��Ț���v��d����x���k��^�(�O��z���	|{��l&]1��۶������vL��U?ل	3Ԅ�q�_�O�p����}GLZ��
�9&w�FM�h��������T��M�vX�Q�����#ӸF��v�?������2����O�Jo�+b�//�Y�{�h~��vgjkA�)�g��Δ4���x~jF�������k�OˍO��v�oH�mh���ϧ�l�XF0nw�������n6�=���d�4���	�;�r��Zc;��tMT'g�V��� ���:y�h��cd��ëɃ8v��G��Jv3���]�0�Z��:Py>��7�`�#90�CB����E�F`t��/�+!듪�Zr`���F\�򹪙��y �2�� ��SX�!�N�i��F�V%pZ���l�����&z�T�:�$�TlJ���|#{F���Ư0����k޽g�oX~���&?�7��_�H���_�cY7
���������֖���$���
�A�bB��XN�L��ڂ"1��^Y���z,�}lT�ڝLS���{q����-�K��@�p� :�*��X饸�����X�k: ��j���!�z+��qT�q�Y�߯W�6�U�oi:����v＼������ �&�?�v�k2g�OT�oj�+ *�#B�>Dr(/��]���N��ʶ%�/s*��C�D6�n7_d[aD|��8+�RD\�:�|�(�O�b00��N�K2�W/��5U���LݮKF4��X��o<꯺OW7� �����ڶ�I�W�T�5�<��S�����T}7��Gu(�^�������(ڨ�[���ap�|�9�h�$�-�0D_�J.����\��T�Rs?�!@q8GG�܌�4Ý��(lـNPx�v;kwXm-���k"�N7<�y�(
h��;�[����n��#���A���8�{E��/�� �m ��\`C�<>�E�|7���n��@�NU�n6rEJ��d���A�HY�m�4��fhjI�H�_�5���	G�;Ym˿����X?��6�3������bY������������'.�V�6O�ҥ=�}�^�JH�xᢩ��`���;�/r�~:} �SȀ�ϓ����Dz`Kv��䉈5� ��1������h�qs�Gk��L1c��HZ��g���y^v�Қ���hW�I�"��|0}�i�&D7�f���mcF��
Ǎ�Ѧ����_R�����_�O��􁦁�І�n*o��V��1�6F�-Z���|-(��[D���L�h�۞4��_�e�&�-�
,/}�_�юTk�S�V���ϟ?yHR�碣\>��ʛ�R �9�q���u��+���&� ]����5窟=|+;��O��-�b��^\����/'P3�����ܫ%��gBl�Q[����f'P�[R����ۃ8�d�����tl0O�1<�X"��Ү�䒭�&�\�A�7����T!��k�tu}��bs��X$�(\t1�n���E�s?)(/NV�9+�B}-~�'�ѽOr�]&U[���#�7Ԓml>^�-�1R�l\�_�G� &���m�ņ�������������R���E_i�0z��t�=
�j��.��m���@C��>?\թMĭw	(.Uy�M�W#������&ؾ櫧l���e����T���bU�l��q3�}�������3=8���L�z�����7�����/}5-h�����R�i7��dQ�`��~�C������������)
෭x���!���V����T�ƶև]�/�c���cԏ%�W��!d�,������`P��֬�#Z�Y*�]>33�B_��o,���5��v6ڸ���p��顅hҧ��a�h��ĩx�Rn�ê�|:�*�'�]
|ҿ���#e�Β����9�����V��s���k)c�����`$��M���Ud��ԇ����e�93�m^I�S(i��AS�V��������Lp3�����.���K�6B���ݹ���M�D���
�'��LՀk��7Am2�3�Y���f~�����{\?��@;���ίL��q��b�/��
/y�Z}h_} l'�	�u���Jxrg��<,yp-Çu�
��9J�!�����8��R��l)(++�]�Tt9@�1+ta+#������ M��__37J*,5�pm!W�� ��M�O���٩qppBm��2�������5|��a�2Q���.��/Ʈ��8��U-��̓��Uy�l7o5�j#y{�
�׽�]8C[��B}6踟mN%�"�����f�8A�S�#��iQ��0V�aק9�jD`5�ȯW� ۜ��,�F\�r����t$0�1c�dKf��g�B�߾$��o������T�<�G{ş��`���!��|;\�������-Z�?�m����`H~�`}�7�nz�`C�C�޾�U����7.1aww�H�~� �]\I]"V`j��5�f
U7I(��q�ߗ���|ىI`=��X��7]FcD�pP�6`f�4��β��ڊ|�j�g��]�хe&�Ω���6(�w$�I�W`��g�T��]�
c�3ۭo��߻��E��GTt�x�hyi��#c��f%�;o9�2E��GO�^�^��Q����h�e�YSUvu��d�������'W�)m*T���
f�\�<�?1�]ï��곺m��R���ߑ���"����T\�vk�Ό�L}N҄��Ϛ�5W�\*���g��Ъ�P��ofsp�K���b��~ŋ��B�Al���x�H&���?̹����zv#�as+�����Xl��Ƞ�L�fl���	&f����;����_m����+j�U\��z.r���냊t{��Q�ūJZ��l�2ޙ{�*K0��N��c�o2�F������î�����}�ΌR��ښ�>���O~��i�F-u��d��s;_�i�*7����0m�W�(3-�vP!R}�:�'��];�D����|�I�*Iq�K��W�E�!?��6��v�FZ��m,��E�2�[���8H��&�!��}O���S+��W��G�S\����U��VHi����_��X� p7�(6ല.�2�m������4�������1�K^���ʒVf~y�I�"u ��D=\���.��+%� Ga;�^��r*��Ҿ�'���s���u�oc�J�J�ugO���Ě�J�����np+�oDs���lw��+��PK�+�C�8���hx�� g��d�)�{pD��_Ƙ�0'�)�z��R�J�%%{�|e+8���6ǿ�m��d��=���/����L���> [���N�!�C/������/ӫ�=��36�h�r���w��ǽ���s�s��|Br7>�u�B�!.)�	�ڟ�P�P;����Q�n6�{�(x��a< �-��W���}�3\�۫���H1��|�̚eN
�	Z�m��'v6g��K`�3��l���/q���ޟ�����/4'�䱥��E����d���N�a��hs�L��U�H��p�ĤQ�vx������Z��^�ÂF���~�]�RLa�_4�!�埣'��?��sO�)�4,�����ܪR�h	+��o���z5��{DG��0�[�vG_��7j[�E�����0�V�������L�Ay�����ư��c7K�&�OHg-�}�}i����-�v�[Y��Q�e5bt��e���6n�3����`�ӫ2�����ޡ���5�T���Ǆv���%?Un5i��҂��3��x��x��˞(-��Պb5���q��Al�O~�ٟ�g����^~��!�3*��n���z�ȯm�P��O��}�l�x�뾯�[�5m��V��Uq6P.9:�/�w�3R*S��ll� 9���芆�ш����Ko���C
���`E���g������i��è�X�!����TN�op{2W-�ln%_Y�<�.6�81/�����r�W[OI'.�?
?���`ri]@*��Tf޷��vf�cq:��2�N%��r�O/`�s`~��C����(�BvS�1�k�3҉����V4����n�96}�y��#h��<���`m�MO������1�|n���G�4Լ���/5��-�V�%g�p�(���q�����}�3��^����*Ї���vcqu��7ω�s���^՟}�o$K���o��˖��y�����4tFP���A\5a�o�>���K�h`�z%���l�=f ��|�f�l��P��v��Q�P�:
�t�xL���&&SI��C��f�ܛ�g�]ޘ������r8�`%/���,��?�@�ݪ)�U�@<"ou�����|�Հ9c�G��L�ʒ��{�UA3�U%��9����E�d������;q���[�Q����")B)�P����[����<3������}Ve���H��+���m�=�Cr��Q����t�Z1�����5	S��2�u�R����]5���<��l.<(���ؙ�r􃇯j��'�s�^���f���5����΃������5r����y�6�yo	.��O�o����' vEﮍ A�I�|f�+���L�I�ir�P����/�cu��5��<�զ_�8+%;��k�8m�j.��ԇs�%gDzF�v��}�����~U�.U���w`�b�MJ���9��#"�j|VsC?j�'Oph��#d��OZ�k��~���"F�z�I��nO�Cay}� eS������w���܋�af�h����mr�^�k^�͡ߣ'�ȵ���E��%+r�~ߘ�GM��t�E�CX�̫�s73	�G-.N2Đ���f]L�Gb�J��7A�K{�3��ށ6V��_�=Z=�"6��Y����y��ޓ@"����de\V:����	F]�V?��VVm�==�����χɅ�x� r��mqō�p���g?��7��f���x�W@E��4�QRIW��<d��s��������sf.'\�m<�I`X���d�7h�u�ݲ�Џ��7mϵ���d�tD�y��B@�� ��UB���̪��x��鮴M̧�+5-?�WӰZ���z�/^+ ��'�=Ό��~��wk0C�Rׇ��]%����a��/̎6}v�}��
�r5 �Lp���;t\���1�V�����)V�����:�B�fS��G�� ���1��\1�gZ�^�X�i��.D���۰���d{s��7��3���O�S<�4�|I��(�NiwV�N�5\�ڹA�{έ���x+����p�?�0�,P��ă��Wv�'2��rY���&�#��!ئ����7�-����R��Y7�m�!U����Bx��H[��M"�E�X�6��v4�vd��+J__O�`]�ycf[9���<XM��GӰ0�#���B�_A-�EE5��������K����#�P��qo��/X�]��f3��Y0;�r#DG��B�8в��� ��n=�e`�7�}�����8��L#[r�Y�y"V?��'��Ȓ�� Ő)�L��&��#�p�*�\�<	-s��z�lN#����]���
���Dч��Dpn�О��N晧`Օ��>|ժ�0^�T�
�Re����	;��I��Tl&�9���KQ�!��.�@I3&ؖ�Z�6�MÍgexq3h�MI�y��Y���u�?oc^k����X��8���˝�m����Y!�fW����>Iv�< Oé%K�_����*��5k��ޗ|�TQ@9MAa'f(������O�_FuY��i؋�'l��f9/�M-��E|�) %0����7�%�^&{��#Ԧ�"��*\?~��0{D��Ʊ�+T��J�]n^/P����������a	��;2��A?@sqg�w}���E\΃�tb�q3��ң��� �W�_�K�	�)v���g�<�O��kX��ޞ{��H���lK)!�A1`΃��%�~b��a�r(�#{d�A��vNw=>	iJY��6[r��0y�Z��36��� �0�r�K`�����n��ER���j�^�p�<��0�6�N|�y��tE/E���,-}����i���N�e߅�^��7��}�2Jp�mM�[��\B-�< ؘᩫ�%ѹ0��uދ�W~���f�n��NDǭWy���2wGl� �U,��ݍ��S�"���P��E���cp�����23(�p�j�꟦�ʹrɛL��rƭ���-ȦR!���[H��t����~�ăS] �`�@��[�-�k�B��.��X��&�x񸽃`[��{e|m@��p��vaO1�Q��h�w)0��{ҕ�N@g��pY_�{�qY���S�����hn\E�h}�>��;��˖U�/^���M���9N��&�O��:�/�N�L׵�4V����|��\㬂��:h'����C��hxcvT�ߋ���
��2�D�&��,�w&Q�Fv���-�V�a�����;�0�?��X�ͫ�^$'Q!��K�ׯ����9lM�LzdI(3G�dv�V�P��̝X�K�so�/��!l�N�5����"h�9����&2����JNS��Y!K�����r���?Ձ<�>��H�����piA��k�9��i����>����e^6z"]�,�|�o��n (��ڏ�?�=��Ӳ���|eU���[�ᴙ��@9����܅��'G�`w�����Q-�\D�{�m���ْk�5]���#X�ԍKϠ� O�y�vl�R��3�>k�u~�>�%w)��k��~���:��UϖW��\><��1����2,�fWR��Ө�����#�s�� /��*ʯ�x���hsa�F�l�(Hĥ����H���?��s��DKߪ�a�W�[툣�����%Z�,|R	�����ƚ}�(������a��i�JL'�<�G�Db�k�~W�Ί���e��۾�زQ�0WȻe~)D5�+˰�Gx�E]�,4���b�˟`r�����g�b)J����|ޛ8�%s�ecY��φ�\��Y%r�>�ݯXyZ����7�n,�6�ᕐ���������ReE-	%f��ok�f}�V'��M�j�M!{c�J���Wj��rKh�����߬�`�����"j�/?��9���韺k�k
�<��/��ݡ��[~��M_#��K?Xy��X��D|����.����>@����aB��9�E�Yx"kK�t�P�#oJq ��'�<�72O[ ��};�����Ȁ��o׬��ՙ���F��?��u�P-��ǟ�0����U���r�����)0$����9ք���-���5�4Y=�F��p���7
`�j��4Vz�e|��m�.�U|�ʺ��i�M�)�H�{O�"�]F�9�˺�,��:�%T,�;���:�`�p++��#ĬC�%�P�?�L��q���7�, >��?KɵwJF�G�������Fy�G*7����=�����粌�l���G����T��sF��3�����W���a �W���|!�)�֍�g7��#8�ۖ���'����Yo�<=}�>���$��T_n�'�憠;������~~���+e19-�?X�a�'�/�W����������	��-Fv�ۋ\ъU@��g�5'���U��2L*y��Q��fk=�R�n�VKadH��$��<�X�K�^(^�{TN�l�O�Yo�i(�l�=[ƭJ1��/����A�<k��!���wg�Z\� W�[�=2����ӓ��3������%.z�xx��w/J�K����9��Hמ��/+��	T��,�Ҿ�-I�{��e��ͨ�L�znB�W�(��ʺ����<@X)�^���ʉ�]̹���x��.�L��X�LtQ�R��������3�u�MI5iX/��uZ��V��6��u�U��s�$4�e�$��`p�����9��\��J��DQ����0)?(�	�dw؎a�<pU=��?�b|�V
�37�djߟs`|��#鞷#iwa;���ndG�P���z���x���zuV�BT�bu�T'�g�@L��$j'�"/����X`�L���)>�5{��Rv�#j;�ztΡ*��b(F���K��b%=.��T��Z�L���S�b����w:[/�w����d�6e:�׉����R�B�9��<IA����~�AgA�:¯8�/<�͉T�!]�hz���^�8L#ll�m�§+~�(,�:`�.>��@�\R��U�V�O|�-�y�d�=)�B�.q�ȹ���[�A���H��Rҽ;@�q|� ����n��x���� n�Xk�_�-��u킝��N�A�rw�\ �/��敏_u��e7#}`)���-+����@������$#�ԕ��,<�����'Tߕw���u��k:���}�����\�}8�0Ll�@�"�a���a�1�����嫧���&����u���mI4���G�Sˬ�鏓~y��"r���=|ex��������?>|n�ݤ
�OwM�lb��'��x1�.�;Uѐy{�	m�bC��S�-3\H����TιD�}/:�+�/���T�WvEڞ&�����Ν�e$2|�����M���t���ʺXC�r���.�\���<SVaɇ��YO�,˙D�*��}��q%'l�ږhR�F�80�a���q*s�t�G�yٍ�$��N%�Pw����A��7�����z`H�QJ|�ك�oSWiC�Iw0�-O��L<<�z/����3�}��hAJ��
\_ܮ33�1"��!Z�a�T���;����0d�ZY�����3�.s��G�(���ط��j�m���:s�P�MG����d&p:�u��WedM���f簎����U��裍�����b}f�}s�m�ٷx݈������5ՙ&�yL8M#���8�������Sq�8�P��w^,ߕk�XM�I�tW��
K�as�����y��QG
��Nt��pȤ7ޖy��Q�l%Q�l�Ÿ�=E]X��sfx�k#l�݈,�p�;m�@��KN�0�2�Pl�U��h	��������\��x�6s�H��M|���r��0S ��B�����Yٸ�d�ct�<����gK�z�����1��H�aK=�����"�����L�@^��v�ZZc�(��MM�j=�0�mÝx�>���� r����K��^V�u^� H ��J�r��
���W�����7�x����P��5�[����7f���#W�vqia�ɡ-R�Q6����#���Ѝ۝�M�w�b{�%���v�f�k�dq��[x����׈J�e�����>##&�����"k�ŵ�*OU�}�P�lcX�!'��Pw�B��G=FK��xCh�2�m��N	��T��b��?�-g�R#�-$�l<`Pz�d��<�W��Fܸ�'�#+e�6�-i$d�[�<	�w�sA���2����|, �ѷ����
1L�s���-o���0��	�^8�TƆ���[KQ�-n/_}"FHGĄ�I�-}x�՟���	N�f)6I�	::"�=�j��;���t�:h�\J��3��\PJ�mSU���O{�z
d�T��C�+'-NZ������:��r�Dy�H5���x��M�{Љ�D���Ͻ�5g�>~,�\���$��%�IO�P�sw��b曲���Q���c��PE��p�@pel�#�&D�1:��*���a�wQ��Lm�sH������Z�!����X{�M�JngE�����`*,�8����yw�c�VrC���;���bE9X��#i̴�x�?,C��	�$X;L�~0��RL��m����=�c�J�	^}�����@�� ]f���@s���o����Q�Ys��V.���R���������]x�ω�;�B�R,\�H��|��}ʱ�q�>D/܂�u�1GXJ�4�"��d�*�~=�Q`C;a�z��7���~0..[�v�ƻ_�P�PRR�sK�j�M����	�M���^[�J�) A��������I%Ay�M#~��Y�pIY�p:j�̗�<׻����#�B�W�^�������ٜ�~�zG^E��ad1"��O6�cv�L��ަ��"Y!-�WT������+4��%|쾘�}�wu���]��D&���V����1fDǷS�{6�����b��J.�����1������nQ��y ز�J���`�bЍ��?�;�>1r'3�i�	�4����Q�Mw?G��7)�)��@B�+EEyT�%K��D]�,)j��%Z,D��*��\k>]�� G�6��1�TČ#	��f<1���5+)�V]]�on�(o.�QQb]��J_gק_3��|�8�Ɇq���$�?Q��4�Q)�}��(���=��^j���]0�IY>���}D�K��b��%4���M���|4�V�~t�̾yh?�����:�|e�q�z��R��e���(imi�������Z<y��	�%���n�Rk�z��C���r�
:̵~��yz�c�gӺ|�ϙ��
�2㟐!�����X����%�ѝ���:���6{7��o�ם�oU$�yƚ�e��Q�r�N���9%�&�@y�kI߃F����R�_A�Ɲ^Y.���;X�P��s�_c�]k���EU��!'�u��م �I2�T�&i��TWJ���X�Q}��o=<�:�i��8�+Ԕ�����"Q��Б�z�׻��﫿���Q{��t���:Z�ʤ\��r�����^x=�.'���D�ޅI�+��8@���ٺ�^m�b�ӝް�%�V��]�^�s����Z���g��ßN@/��� ������W��؅�c4�!p�.���fk���UH=�=����y��jM�ȹ�::{���r+��r�����IIz�M�Ka��|��FP��D�g���ЎMn&LՃ�����o�\R��zY���c��GvI|D�.d_KV:��]����g�	�ʱ�
;��e\�s�8�<sΖ����#)%8H��U�~Okb��9�'С���1E�Iĩ����^0j�_F���m�=��z�yrMe]��s��1����SW�a�
@x�U{'�������28OIbd.�;��G:�PчJ��,'p�5'�����.�6p����̠y&�� ���lO]��C9��Ek����{�H2�:�]>�pj*�"�[�r!�#��0�=�9����9ntͷ�}[7��m�8�3�k��c�=�_r�Au�{�~'S&��WLP,렷�d?�L��9���$�Z�eA������5'��pt��s��u�Cd)�C{��DH4}ھ�gHʕї�H�{SE��Ʊ�����WL�*��ϼOC�X�����pW�pl���b'�厌Kt����:��O�v-�������?�Pj����a�6�dKM4b�@��ӿ����b�|@���V�NqӵD�>�12V#`�;Os�ߦ�zI ��5T}��=;{e������E /�`�jV.>S����(n
���_�<%t�=�)]_�)������w�p�ԇ�{+�~5��M�vh?��l��/�ŋbh�5R�?!>X>'��[�v^�����u%z���;�,�Lu0�g�@�;~�ϩ凄��&�w�te��r9��z{�*I*{����!bν]@�(招�����a8��[�Sp�Q�d�=��o��`>������e>y;N�z�R3q>|�����~)�Y!q��n����E�,(���&;j� ��~��E���m2����5�|�&M���+r �W���]�J�)��=^I��8l]���˺����ѡP���1�3uD�$�KL�O���$wd
q*����1���ꆈ��������(�p�RR?�!�F��G������('��O�$ߒZu��{�6�iY�����6R
��ft�I_�� �>�mi��Ԙ�����Eu�A����ȋ!.�[��N�W#�#�et�?I:p��T��Ӿ 8�Co�i��6�}-�O�?gf�SRBOo?��5���6��7ԍ�I� ��}���;WM��D%L��LU�8��U�
��<Ȍ�T�^v��(��#=o�*�-���S�"^IY �1�Ig�
�Y^>�}�в>`{�O� I�&�t^%+�G�~×.�P}a\�r�ے�\wmc ��yN���z)�n=�&2/3�,�����Ɏ��ر�G)}�;�����V:!E��}����u��e��hF�t�9�g��*����>O᧥��k�]{Y���b� Kh��A��v���Ğ
~�:�ړ��:*�%�0����gRG�+u$��W��VT�[-�
:lD�=�>_r��Y����Y<IR}�Ӵ�Ra�e:��<Q��� ��ZN�}=�}҅�	��0K���Ug親8x6h��3���?�W�kV���	���Q���W�S�,��Va#�L�Ie�@�'�3�D�&;�;{7�޸G���~�Ho�_���q2q����K�v��-�*|y����E�f�1d�������^y��Uf���,���/q_����d?���+�����
0�F:�[�O��oso�����>)���nڹ��@y~��<i%�+��4�U��(��q��\�U_ ;_6ߋ�\��E�6?��Xg���͠A7�$i�ޞ �ZA!v3���||օǚ�WH8pJAn	}�z=�tX�{�q��TY^Y).��<�'I�6��z�E[H��M^;I�7W����yKZ*_��@8�+�����7W�,kj��]�B^�,�o�s�4�K��3%ջ�:��.���X�Sv��6}��?����#�-�g���K���/Y_��}��PVZ*LS����>��z�r�۷��Z��o�wہMj̍����TV|FXN��E��ӥ?8�j{Ŧ]���C7�K]����N_N�P~I8�K����K�R���/���O��e.Հ�SWK찥C��b�ɽ����tqth�.�i�o6`[��~8�ߓ��q0�'$�������̗���
/��i���$�-8�\� w�_�����奡	��Ѯx�?�.}g+l�@�=�=p����ZX��V���Yb$=2ݩ���^�dT,�ɼ�ۜQ�]�<^�{�.�q���o˵T�v9�����)3���i�Jz���3ww�����l�%����iz=w2G���ʟs�j���x}!�{��h�]�	�%%���FFF��=�<V�C��?'+DR�9�؞~\��*�����
"��/(�H1���&{�&��0=���W5=�59c�ʮ���]z�m�L�˳&�}^�����<Yd]������E[��Lt�L��z"`�r�<���>�zeU��Q (!�f	ڢk�.K-x)�T~��8�fo�^�e�?6�M��R+1�c+Tcb;�Α�g����E��������⧘���� �*r�dr`@�:+�[�ǖ�#s;��p��<L�	9�me���_�q���E~�������#���U�<����,~k���R��;����S&�Τ��w�K��4��޽̓���*������@@��w���q��E,�����O�5��co�5$S/n�Фy�/'8^�-T�/�N�]����r�fl����G��+|4w�s���u�a��y�+$���M�pw�LF�����GY�Y��c���C�'�������ր��%]|||&Mhd�鶡�@.tn!Z�%[�o���h?��/w���hO�G�xڲƾ��V��i^�s<R}kC�Ջ��F[k�^�I"qO�Ύ�pb%lt�")����V���N*��C0��uJGo�[�C�y�-U�ևYbC���R�<�q倅'�E��,�Vb�Ј�΅��uI��f�!��8�w��;ſ1�lY	�=C���2�RÓYh\����6*���>�LG���14麇Pc��Vk'�y7�JI��v�C�H�+���/��S�xg��2��dq��,O�H��d��(V���7شN��oF�L����r�R)�:)���1��܈2f�A�=�(e|�#���$�Z������M��w�A7��9��#�K� !�o�A�=�f�|�+6��\�jI/=���aC�#�R�ԅf�>C-�x2X`���]�)�x&f�c��A�f��P�aF����%�G���d2���Aƕ� .�9���0��0�[��O�W8��8�Qk�u�H�ċK�b'��~�x�V	d��	�8��O�%����CŻ�����Zu��?&��X9:Ԫ�&�E	���V}뾉+,k	�by��u�c(��6���N�mI�-���ILYX�!h���e�������c�y��u����_���!�0ic�B4�I�Ξ	~�a�X=[.�8��nO!�U�I�r��[�b	���Ѷ���_Ðȧ�<7����k��V�s���l���W�Į6%vYu�FB6%=� P��cs�qc�ю�ߣ��ƌ�c� 	;c�+�[�X�E��;ӑձ~bw@���~�u4�r���[�z�ue:������z�<)fM���-���d���H���CCk������' �z���B�r��jC!]]G�O�h�*λ���5/�7*S������#���|�u����Z�{=��o#@b�V���>�
"���mg�;�$�]�ײ�����:9�B։�n"DۺS,��Y��^�����G.���"�jW��r��V�L��@0���HD���(�(R�̃�k��ŽF2��7��F�!���^+r�эM.�c���Ճ8chU
�&���7!����+%:�Đж�@\��e���B�ʽ��l'��D��;F؄"���M�o��"�B`7>Z8E+]9(�b�ËE��f#E����5\2�x�V1����P�H/�,E�^r@B��̆���q�=��h=�J��[���Uce�5+X�Ɏ�%��
��Tyܖ��9�'5�����k/�8��L���e��W��9P=�픅��o�h=G�݅`����v^�l��Ţ�.&�̈́��&��f+4A"w����daU4�Fv'�"����d�_K���[rPȴ����~�g��7�Q{��2���k2��5�(@s�ܠ(4З�O�a?N^���k.��#"��g!cr�����?��x�{���JӶ���M��Z�����+H=���hs����|Uނ ��d]�(X���Ϧ�;�O<V"n��}^`_USEdFh���Wj�Y4���5H�K/8N2�{��)�߯��$�4�4�0th�4��n6p`�K)��-�R����Hԓ�q�ՙI�����c�G��^�/PK   ���X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   C��X��iP  K  /   images/e6075517-c690-4ca2-aabd-cadc5d2d7233.pngK��PNG

   IHDR   d   -   X���   	pHYs  0�  0�
�D   tEXtSoftware www.inkscape.org��<  �IDATx��\il\���6���vlǎ�8���',!��&*��@�JCKQ��O[Z�U%ğ��P���DE�P�hÒ&B��4�N�I��3�Y޻=羱�f�č3�`�|�yw��;�{o��?�O G�鉿��T
�,F��I��PY�Àl�r�|*G�T G٠f*+���`�0 T�T�S� G٢a���1ѐZؚ�R$P��"�P�UL�ꨄ�Tq���2K�S5xB�Pc�1��������d&�6
�QTw�3�	��,�dDE1��(b1W�:S����>��ē׉7�T�/4��cě�1�/�|�P,s��I�&����tł���;_�2�G�h��
�x�I�A�-�-��ϖf)f�fŊߐ����.��
	�'�<!�<�'H�Du�����~���j��f}�k+z����U`w�
��^��;K��F�ŝ�0B4 ��¾.���Z4��G?ҖtC����׆��D���i�Y�e�6�/������ð�1T������#G�G�0�Hנ�# ӔԮo�oG��7a�{:�T:�����9��$��M���^�m
{�~���b@�����<0�'�r	������n,�����7�;�ݍ?��"��9:X�R1� Me�.�,�R ����!}!*��^W5zB^�RB`�r���\NQr���&�6��/�'�}�u5\�c^D�t7#��P`zˡ�%4����p̣�'�2t���N���f#2qR_'�ƛol�S�«����;L�䍚(�h��O�1u�T�r��x n�2bK����n2NO�)��2��]']��+���Ε�R��۴2Ϳ-�L����g�h�#�L3n/GU��x[����oa�2|�[����ϛ�ġ�.�G����f�nX<f��,�_�W�=�[����:
�c%��H�e���U��TE�X�p�6���J��*mD�~V�\2is�9���ϨQN�{��YΥ*r~����Y�Te��(����/�C^	��*���+�cPw�SY��/އ�Ʒs|��b/\��1��7��i/������s蚂�ZD}MttP�[p�#>��b�1n��iS��Q":gN1����l<FLT�j(*�ʃ����6d�����R9��I�zq�m5x�߇�5�`(+	H���?h���܃=WH�SR"K�wei@2{ Ew��������4��� �z�r��X�\�7��P��0�yI��O��`��q�K�k��5�m�q�kv�<��y~7ml���-m�#��,�p�����C���Ç"q,_R���81��儬��]W"5�rv�$�Զ��#R�>w.�)Ǳd���@`���y�ĸw6Ǒ�N���;�"�i�j�a��*�plk��{Z�|N9VR���M��ה��d!���i�o�l[�5�#w��3q��P|��S|���j��q=fNϧy�q�
+V�����w�p6%�:3:
�*��2�\:0x���{��T���b|��7no��7J��(�ó�j%�_x}���������5���kh����^��Ϟ�%�K0��.�b෯���kPR��/_�T2��u˨P5ݏ��y���_?s�y'��:�޿ �y�Uy�,<��:y�x\H�[{���B<z�<� �Z���5���)~<r�\<��6EmA�uI�V����?}�F���;N�3o���kN�@[� ��L���������@�l��%�Ȕ 
)��gL��<�����:p5������+���#g���)m]�CXD>b��)���b�Ԧ�E`������jƬ��6�؟���PT�o!�h�$3�v_ɇ�uؤ����y�/ _9%@��'�g�`�_`�+��m�m�h~c�4n	ǂ+�IA	�f��ɹ�'������4�l	&#>Ի,��;�U��`�������#+�N�aӮ��bS�rY1�;?o��p������X�7F ��i���s��;�Y�!��,�a�t�!�6v�d�?^{����v�[ 	��m�l%�G����	��\+��mn�>�l��a�	t������X�t���Zۃ��Y+%%8,�z����K����&d2��I��dY�Q�r��#ܾ����M�>d0��Zq����F�������
�USf��PU^ �v��Vɤۮ��~�$�@>0;K6Q'[���T��+����hEiQ@FzX�I�(��Qo���7�������E�����?Տy�S0��X����
S$���F�?�&�d������X!�VO`��FuyiR�<#�)���C~� ��}���c2 P/�	e{���[���H��B;oH���Jں�d4�S�H<ž#�h8�Ѓ��ݲ�c��e�鑼C��l������Q�x������Kec+�h�R6�9�&�Y��퐟9l1�O�qlj>�3����#s�>�&�ە�#J�f��&{�j�;�5������;�G6�{��zEu�T�����L�'2ַöQ�Re~b�T�R�i�pD�v��4�2�0e>!%M�y��X��8�?��LeI���
�/�F���1�t���s��˴} }J�*ι8*��T�g�?(:_�8 9����2� ��D�r���I�(V����
{6�ux�8�3d�o�y��1�e
ѴH?�w�CKd�|-�Ɣ>�Χ���G�J��s9�\���q�1u��2�Zv�g�I7SL�2N�<�};�b??��g�9�d<I�'O�����sL|>�_P��0ׅ�)M���=# %hZ��6�3���/�D$����SNӻ����my�4b�]tůfN��o&���P�%�����i�g����х���-MF@"�H�E�M��K~�7m{�@�Ӟ���|��CCCC���ԷN������P��U����N�1��I�E����n�1��þ��<&^#她Q@(11]~�-}�w�HA����^T�R�0�%E�4Û���3�C��k�����dc�]5��FKsy�/���ϓ��V`��� qß���`nN����?�%!/��W���DZ�d<���>*%p��'Z,�C��=&�]!�qw���P.���<A#��w�G=Jr��F}��o��xBؙ����1/:8s���:Ge�԰(T�gpyЊD�� j�?�Q	�E�	�[=�|1�*w$*�a�r���q�V*�PY29i|D�.1��烰�y�������r��e��"�f0��bv���KAK����r��``Y    IEND�B`�PK   ��X�3S�u� �� /   images/ec43f2b3-9126-4f13-83de-62ba1ea97088.png,[ct�]ӎm�'N�F�ݜ4v��m۶m4hl۶yb'_��ߏ{�Z{���5��v���wd000d���"�5�!��/��!�oP��e����b�������Jj8��������P��>?�b�ʮ��n��#4��U�/�::ͭE���B������`�B� ��H��ia=�O��]-��SA>�r���h$�P���`�&<8rvIr�/U�eE��ww���*��˓�N>�rk��r�/��-5��G�|�n4�u?t�о�c����,���vBɽ�]�8����o�ڸ�Ot뱨�ڸ���O���k�zݺ}��P��w	ʃ}V}��}b�?εf��
n�0^l��}��xC_���I�Bȥtb׈�)"<�~z\/C��伭ɕ��/�Ĭ���.�-m13ȕ=]}��y�����}`�}4���z����c���WR��v���fo?G�A�-E�[�E ��!����РQ�|���}�H��#��"����7:�IONC��������j:��cI��U�g��oaŋ@���H���X��Q�l�_p��&rZp�6Z���;��zh4�R}HM�-�Rz٬!�7�,��:ҠH_Fx����r܏M�ȃ���i�
��������7&3#�$p��5���t�Ҽ��we3G���
Ǜ!ie���XN��o7���c�D+f��#Gߓ�[��#�Q7��0�/V<	,�5�+���w?U�J'1���S��(4#��BVma3�.��{���]�(c"����j��Pg�3d�C���L��͒#�����_	_j�?wG����+�z�C�V�D�^b��עd@��O��-�u���.�9�+�����U~"/�?bš0�`ꦇof�/��\zc%�_l毳vSG���興6g�Vq$w�����8wX6J���2�1���P�&w�߅Y�Wz�	���l�)������_Өƨ�W&�v����L� �\bK��3[�&��}f3Ls<�S'j�6D=c@��m�� c������JE�B�&_{�����MB�x?��Cn���s	r���1�JB7��Lb��vuś��3T�"�A��|��Ee(�Ϟ���Δ�=�����d���U.��R�������e!��k��~���aQl���<��B�՟�K��Ɣ����g9��.��=9�i����A�Ϋ��yH;�N�YX��V��)>��ͮ�f�%Z���[���_�"���h���|6l��puȨ�}%J�E߯9#d�FZ]��W4��� �����>��3Q��5�E{f��ylM�'h#�hFPֹ-��=v��˔��6`�0���f��g�Z�41ȶ����PC�+����'V�HG�|ք��CG��/�R市�Ǥe=��?կRz�����~�G�>�0�%>�w���i"z� -7g"m�p�Et��`m�hB����OW]$��۶�p��n}J3��D�H�~<���~Ȩ�����mY}Z7��{m���x���s��<>_�l~��[RؚizKE��0�G_[�?N`��B览c".Z�YU��n=�}xj}��8����_	ތ�y�\�V�۵!߻#��&D@���I��T��������υ��kР@���6�M��އ�������6�+��A���*����Ԃ��ލ�Z���#�06�t�j�!���ll��ԃ�}/�����t���T#�%&�����_Q���Q���4貾�g�����y�9՗�ۉ�x.#a>=��n��حY!̰d҂�vuѽ�6y����F��Q0��8��Q�_�
���]@iE_g~�5�潆���?��G-q��x��-�����1�6Y�\<l���<x�Sg�q��F���{������ۇ3�gT2��HJ�x��uF�n����	��:7�.r����;�ʈ���V2���o24��
t��r<]���n~��<G�-�w�V �o=ہ�H�Z�ݷ�jϮ>����_�0*^�6��3#r<ml��z�B���Q�A4��Ln3n�8o�6��;A��$���z4u����w�Y�L��\���2K���^���7�	��K�侂DH�9R��}�{�Z<?��{	�5��`k9�w.�[���ۯ��mvUUv3�2U�`F�e��l�������d@�k��Hq�JmS>`��ji�_TY�ᥭu�<���n���9���蚱�L�!s\�K��8�G$fp^�􉹣�s�G�,r�G��n��նi��e-N�}�I\��ris6��m�h��|����Co�}���x_��0��Y+����Ǖ��!��*�(rB]���jM��r켠��E��cs�E0���,��U�W�:$w���5���`R�teh�U���i�����G{��h;���Q�ӳ�Eꦺv���O����_w�O�r{����l�qɡ\�!B:a�3S���������)���ʳ��c�j��e{��BM�f?���)	�$P��H-���Vۭ�X���oe;���䌭J��^���sԶ��cK��џ��;n���;3��9�[u��~��e;W|Ԕ~��XG���>_��k��~(�H��E~\�n��[��2�(���|EM}WC�b�����]�IR�4$y���"�s$j��s1&]�����,bV�=�0!9���_��(���z9��iN�=� T�zd�0hB����ק����2�]v�S��'�#:/�;f r���Q�����H�e�EmҔ->n��	�壡��+�_��$����߁��R����l����㔿�l��G�@|
���;���4.��5��T��b~�{�9��cʩ�	�ШGzؑ�̭���_�7\v׋�S������G�ǈ�S�S��+e����[�e@�F �Y�� ��1�]�թ��|k
Zy�}��潄��Eݫ6]�.&_���hĴ�w9�|Pm�>Et�;���	�O��EǽYH�KEh�K]���Jiz�]>'�9�T�IG��?6>�#�9�h�u�)"*��Weш�gP囌63�8VB��+��p�(��q����C&aoৗ�'?�` �2e���-?;0��%���ں{�Rg0|��w(�y�
\N���X}�=����R�V�l%�eiN�͋n�#j�� ���N�<jCo���{��-=�$oR�|�Q�_D�[��oL�^K�L-�5�[4|]V�Q��V��kV˫�c�`�i/�_���B�X[*6 ��F{�iv�)����s�lN�	���A3dS�o⊣�3�ü6���}*j�����r�i�#t!�m�eX|�S��ïp�V
�j"���U�"���~�%�����rC�<hH4:,�%dսR2�BSm�1>�f�����A�Y��r@����������{�u�s��V�u~��v2k�xO-��$A��44�x�7پ� }s=mAJ��4���zQ^��`Ż��!��/����K����h1����=��M��#ա�E�%ԅ�Qi��=�{�,d펷n��o�������"������Ax͈�9`(&	�VӄKBVw�]�q?��6����]h1K݉�g�v#��}��
�t#�rZ������'��(�6 [�e��]�#�!��E��%�X�����BgF3���pF����*����-��$��(��Н�KpW�i͑]1L�iם�a�Kr��[�6�@�D���[�Y��+�c�v�k��+��F`:�w��aa����p�mmJ�Ϻ�ٗ��kQR�	��R��������C����A�}�s��|�*>��o]��i����p���;N��%� ���:�A]^��D����Q�^ˌ;dͰ�/ nf&�C
g��n�q�m�0wm��=i��b�E���Ȩ�B2X��@¸��r���+
g�)-u���-���۸;��I�
\{s������wOEC�&��7wF�?t,���Hӭ��2b/�l]��~��zjb֯���eW���0uiKn����
�8��Ow=	:ߴ"�㛡�mTr7@�M��=�����kA���lN�.�q<k��/��l�m��z�%X�g���z��|O��w�����i����F������`;���q�w4��|�#�y��VaݑBҴȰ����x�f�$0�XY\36�!q�V�g�:�Og�I�;�( ,]�Ä����`C��1x�a�}k���a�9��N�uJ�����Ȇ�#���)�Z�ͽ�d �`8=nh�6}�;�h* �j��TF{�t�}jM�Y�����Y�h��2c)`U�`XS��-�,���N��o�17�B\'�u��iWQeA��Sߩ���&��2�;�8$ƒ �Y�*~r���kO�>��F6��._q7[��k��oj����Ò�������(�p|> �y#�Z���jn(A��mnn(��^��?g��{Ɂ]Ycf�\������6�ё	-'�V���:��w�z5
�@"��N�����:��E�"��;ҬU$��^��7�d���5���ְ��LzU�$�q]_�:��b9�\�sD���0Zw��w4��J1�BƖ=��ؐPX[����'~����<=�_��lj9��H���4 �.y0R	0�M�k��Q��?��hzQ�lJ��#�t�>�������#�e�#RU���j?f��.�]�Zl�Ys�'�V����<W���G3���|
J��j���{���[[%V�*�*�<߉���a��e)����`Uϝsw�y�j4�6BvpX��»�9^��*/o�CS�PtUTʔ�5�Z��셜�MS��:�&�.[^ʵ�;Q8\Pw�q���6�YU�>��i)�k���\u6_
���u��S��1S,�([k`��ɦ�z�R�hߌcJ���� ������\[�h8�����C��o!�����1����Y�����P��Q�ߤ;ȴ7���F�(�v�A[YI@�U�#̲.�R���˳��P���)��9N����2x	�x^p򍋿I#g!Ԟ<�6��W�PɟG'\�1 �݉*q���[���2C�o#^	?=�c[�WDJ�*~dr�#wv	�c���*��Z��>�| �Y�'=`�FX����8���}�tו�Pɵ������a�c�YX�r�_�D5�yt���.�b�,c��{�!l��=���\w�����-z���s��F�~������<uAK%��d
/���6_����>�X�O �������A��I�&��V$�f�O�4��nd��3�?V!�܁��ú�J�����7�ל���v��{	S?�(��ƌ�,P�-�Tia��aPW`np�tm�^�� �̎�/�O�W�[6�N����i��:�����Y#G�!�R�~�,:@���B�������Ցnm~k�w(�$��{�,[���#j��'�`��Ѥ�ʋ���^֡E�%p���_�����D?�*ɟܓ=�����(�+|̸3qO����۪����bX�t뛗$vd�U�W�d˽]��!�?�c%K��.?�!"s
�����"��b�{���[hP���ɷ�g�'f��/	����4��\�����z'�����)��%8'��i$LRh��h�w�cH��E���'�_�8�녀8�2��dv&G���n�K��� ���3��������I:�����0s�kѣA�_��v�⤍�ũ�?v
��j+��� �TMf�����<��Ӳv�eN���]������\�fGR1j/H�"�Cc����"���m�i�_3ϫ���o\Â�Z����V"��ڻU�-�D�ބ�iɦ�<c6�8� �� ->#=���0�|���C�iÝ��I=����8y��y�9�hW1��Z����v�~�x�^-���J�����������vZ4b�<��l����c��ǔ����t�ϊ67�'�,�sr��MKU9i0��P��AX��]���	���ၽoD,}�7�X����qe��XouBW������xOmߜ����RT`��1I�jѿN�fy��?���<J瑟�9f�?�h�|0)� ���ഋ���)����x�������SŌC��I�H�KלȈ���]b�^����3��d# nuOozT�cp09�=rB�<���
#���iszOJ6/���!TL�� �Ff�Vmͺ]:Y���+E�ow��Jma���춍��iM����q!an�� [G�B���i���:�é��BE#���5�G���|�<��,ghłu��;DQ�-��lDJ�t�Y��9���麡�U���] �L�s�c!	�s��d�蓛���9
�s�΄u�Zſ<��Z��ӥ)��_3��:Eb�\�W�K�6�B_�g�]i|bm
�YS����mޑ��	e��wb��T��@��鐪�w����=�1]�etk�B��|T�\Q)4�IlJ�%��G��2�Ra_R~uLo�n�ZrC�R.��}�<qϦ���j�P�.f����OUV�X�30T;UQ;�뙹S7PCn�<��_��{��y"�#)�j@L�i�:D�(�b��7LX�Rd��<��婢D��e �VJDwp�U�j���dⰤ	�6gX����E����^;��5�d���E��۩d9f�/.|�iL$v7�>�_����9�%��;j�f�}��F�D�~���U4	^�R�@ڳwM^�c�Bq�h���M˙�l&#[�D���	�g���ε�|�ǭ�l� �OW
��ꃈ�ːĶG��ˀӯ�x ��h@m7�GvV�;�T�l�ѶmH^3hӟ1h?��}�˟�Ɠ��F����F�]%�����<�P�H�D���7���f�I�Uz���#57V@�}tD57ӂ%`=����
��*<�۟B)F>�5	���6O�PZQ��pB�b,��R�����}+�̑���F�◆�Ax4�8l	��+��S��T��m�̑�cd��i���)g��g�v��w3����⁆�i2����`sG���Pi�-�����}K ��B��!�I����Z��$��j��p��?�U�N¥�?1�~�ӵyfad���]�y�i_�<⫈k�$e����[�c� 8HʓK���XN��Y���ۭ,'y�eד��!S\,�`,�]>�J
z]�4�L�:����ˌ�XeAZu��Ǵ�Tˁ�fm�Q��$.QE����g~�����	��t��t�� 5?��o�ַL���"b_8D�Y����8�I�(����M(sw-��:�C�J�э&�,sG�舙�N�������n�R~��g���^��c����7�'���Iߝ�c�#��V�<�F���Vwlr�Ǎ�b�E��b$�?Y�yɛ���۩$��2Jx�7�f
�V�d��#�W�W���/���]�2�ϝW�F���)�p�s�2K�ꍲ��$k�J\m�'ϴ<�(���j�Z�kzH4^������q%Ǟ��j�Κt�[�\ۋ#�Kɉ�{��~W�5��AA�X!;ù�Xt����1\Y%~|��ȃP|ڄx;)L�c��[�3}�\�ލ���E��rM�No��g,��BE7��_�bDǾ,�ZU�%΁r�$�2��<yUpv��Z���viY5���`� o�|��'nE�}�ӄc���|9��E,�D�Ț�/*EtNI���Ӭ���ۉ�4�ԭ"fH��)a�R�cY�(x�?c�t�'�Q���*lfQdg�0݈-`j,�WW[X}��j��Gi�8����8���Ϟb�@��
��,G��ߡ:�)"�R+6��"5�q�#�%V�V��r0 �4F���4q����\ļ`�׍����P'�[��U�%X�o��Ǉ�8�Y��I��e�1d6�����ĥ� ��V����.2�?������w*����Ϲ�8Ie�����	/���O�)��`�*�P(��QY��w�Y`?4X(���w�D?�#x�Z�H�&�B�(�q��3w%�-.�'�����"���r�1~`�]>�+z�D��˳��p�,�&:��$ZrY�8��w�zҀ�h�"���?�4����,�a�Dy�5���<O3Qi��K�5�C�S���"����tO�5�`!��ɕK�&��\yĤ�Ѧv_�0i�hDB��eV����Fo�{v��0�Ƞ���y�˭���,D.�C���XoJ�
���qW�>�SYn�_����`İYH�u.v���L�����s�֜:i��'.D�ŀ�y�I�����x?z*�;�Ѣ�$@��Q����,2���i��$�$��dEJ<�1#��/�����LP@qZ�a���ξ���q��OZ�᫄dS���G�-Y�;挔3��Vrݲ���qw�ӦW�؊���&�
gd?�r
0X�k��S\����響�}��q�z�����W���#�6}��%=�"-e��.Z�Z�����MM�v�~����O�f�+q�8��"K%��ZvO���{���-(	�}cr�D�6��N8���sV�����Zc�7QP�T�5�!�U�����Xos�Se�w��&-�ܡ�)tBQ&1x��GL����Z:bs��r\�a��PI���Qah����pV�Wk�X�\9il�, �&)�U��Z�9_�d�[d�n=��$rU%z`����
xb�G��e�QS��{}��4|%�WEr����DH�.��/d�rW���X�AIk�����	��Y��B���$�˃0�"NQ��?y��wұ�!��y�w���u����NVU�0<�A��,f�����Ϥs��ctuT夙je����:����Сnޏ���ž�n��«��`4�*99Q5�H��d�̪��TRIze'�ݝ���ukh�Rahˊ)�L��~Kv�ɫ�(ˀ��_=�Q��-,��Q�e4���Ls#�	��ci�n1��v����@U#��)�����UPc��:e��{����?�$�!�6�P��ٟOf�!
�q�p��Ks��.6���	�M|@N�*b�$d�#�� �s���N��Jd�g����?݉�t3\�)lJR>I�b���
H\��`������\B�^��9i��%���b����q������b�Ίw�*��4��	V��H����]����x]�R�+�P㍧s!�F�FqH%֫�]�Їq|'�D�}�D�1�J��:+jC+�rF3�)7��]2���k��\������q.�1t�5t�8��jK'�n��oi�5��I����7���xa፡Z��E���l|�rt�&��Ld��&n.��'��Vs��%D-�#�9A�N.L�c���f��zh"�ENq�z�� 6�*m��Ox��]�'����m�p�Ħ���Rq'�x��Y���Tt�h�x-onN��%K9G,\8��������:��ȡv��-q�9�ɦ�=��4������p�Z�[h�]�a>H]�xά��W����v�53�e(�������)�O�(��ˬ2&�����D�����j�G_8B��y�~f/��8�k�UbϿ�4����7ގ�7�Q� v	S?�EP.���I��FxhB�ykn�����JU���X�&���]��r��	�Q�m��T�7�`�3Z���5�	*8i�������dp"�O�{�����/]��1Ri\������o��C�n��T�(7�xvLY��jI��I�OZ+3�'2����	;�K�4����ݿ�6�4%��MVb/����z�0y9QC$�z��%�1���v5L�||e���	o�߷3�~�����&>K�(�d)��JL�m�ieR��=�Z����Qw�
������O�Gë}�\B��#�>$�z��%�F���$M���~f)��N������E�Գ ?2�<Պ���5m�V�~+�����@ ��)"DH�$�X��1�qJ'y��bHa��a(V���Յ,�dz��L�f�
ď�S�EƎ�3�iA6�?go���r�Y�3����"ι #����ge�:�7�J����DH�~�d�����Џ���=��OCu���U����F�F�4�r�����:5����*ْ��7�4 �*.$��}��n�WD)�*ggw^�h����ICCI���:����k��u-M{@��h���w��l�D�,��㤔��0���K��H�Y�,����I��׺�*���]\pQVC���Њ�$c��X����;��� �B�\�_Q*
��w9�%��xR�!:�����/.n�=#���`�d`����G�����/T@`?aC�]�0��t�*`��D�������+r4~EUz6l�^?2���}I��"����*-�'l^]^��e\�^w
�.;�&���s9�}��[[s]J��h�?�H��g��_�} I���ߎ��ptܯ��-�Էr��8��ܓ�X�s��Y_w{�jF UVt��]`9��l>Kg�p�`'���ǲ)M�焞�k�Mq�}rܮW 	~}�sŘ5T�}���	tӨ���sk�����`�|c�b��M��WQ�S� ��ꆙ��{���i�+ "qm��D��@1{Ǎ�a�R�^pjM�ٺ���TU�4�D1�;��r�R�:�y��	��=���/l�n���aі1�u]�Md6�k��{y�kgDO`}�*E΋p�� .8:�������z���xV�r�p�# ����)�M�䭐,����T�k�%U��1�-u}p<m���	�>P�q���C�P��#��K�k�_�W�� ���y�`���L0v��IG��ZxH4o7J���/�8�בYi���H9e�}I�$d�ǟ���A,p;��������0YM�Yx<��_� E}�m[��-Iz;�Ml|^y�>_�@	�/ஏ���/59d'�<�F�+g��p`�/:%A�($��c��p2vE�ͩ�aM˯P@m�+���DK�p&�o8w��mG��;!$��/�C���S��U�']�߈r!T�w�6\�����9��db:�u\?xA~]ײOS�0��D��r^� }Mv��Y�٨^�q�ASi�%"�����"���b�*� ��#�Qَ	�O3�f�G�P�x�y�T��X,Yw^yq�'껢&F7�&�J��~㽷A��h�2b����܁\��EB�5��ݐ����l�}UeS�?k&�A�Z V%�I��D,��R���8>��ts����-�=�qa��S�M�}#�~�����K���܀^[��\2�Qs�A%��g�����-#��'��&=5�ˬdc�К�󭈹����z���G`T���1�0�ºmt3�����D���l�\h�]j���m(g�4�`��lw(����v>ԶW��v��������V�E~/k��So@Im�K��>|��h�? w}.Jَ����I�����@q9��8Ly'��@{pv��̍��W1�����D�-WH�'��֊?�e��*"[��k�l,(�g��EQ�4���P�< u�wB~A�IE�3q�Pz���Z�cqxb�
���M��(>P��n)'إ��c�p˵XӤ`���d�S<�����_mא�P����&'0Ybg4�p٢���5M�k�y{\�d�|È�C��\W��OҬ0��E�+�������.�_�$4�dkG�w�L��vȵ�u�*���Yp�n�'(��]��<&�vV.$<eqo`��+�G�Z�08��t�l�pw�~��0�Ia'��b|�e-|�7��XX�>��}�MI����6$��(�B�cz�?���X��^���UNȒuT����s��J�o�W�	-@w%�g���m�D�Oٜz�Esa�oAh�N�x�.�z9���܁2���%0s��3��l����g��YL��ps��X2Zx��y���P��Z��bJ{y
���A�a�R1�������h�5�͈��k�Qf�Qi�u#�����e��;����*��v�����F#�/��wA��Y^-���)��~��R�;ze�0KV�?�EC�vtÚ�b�{=V֖�MPw?��XU�1�Gj-�S�Y���<�ܖ�}�C�ʔ��7!� ̀�H�:/�Ɲ��eU��
Ǹ�R�/�ɓ8�5:��4FLIt��s�ln�",�r�j�WۂD��DĄ�_²=�q�zoHل�>�,5}����E(��V���V�h�SʺQ�2I�#��@VP�D\x��|\�,7�U��c�i%�@<�Z�4��S�Cߎ��b1�D�+�A(?��(�gÆ�;\�v�p[�5x�j_&���P{U��'���B:�J���o����� vE7%g_Z�?ư?��#W��s�^I-υ��H$��x�|���tްx��tî�I�}>�Q��HX�f*"�����_]S���I�k�l�m���������/(�h\5򔫙E�W+�I~fE|'9��M�ˌ�xP�0�ݥ2�m=[�\y���ZH�X� ٰ}}�
��M��h8Z*�{�5y����J	�MJW����<4r<�º&������D�lnD���0sNLdaT<�H�mT:l<�"���/��E�s�v�"�]V��\Z�
�tߌS�]8������l����J^�������ob���M�Mئ�UG�0��/ڰ>r�m&�S��Yy�`s��d�/ܿ-�¥���8��P��|�UZ�n���Ӛ��V��>lW�:��˶�'*Ep6���场^<|ˆ ͮ�5ЃKg@���e�o\�(�;6f�`�l�U\	w܏榐��2��3�|#k�_�rιD۵E��L<��1]#Rehvp��׫�Y[����J��;
�XJ2����#���B�N�&��4�'7x��ٽ�V2�9�B��Y��m��Cύ���8�d׿N�~�0@x���$�o�q8*�背�%�NjB�Q��%�H���/��{ڮs`�E��X@��w���*�W���sNs���u���xl�[/�����(�����~���V}h$�N�*]���.R�JH��ȮD�]v���Oo����YA__<%k�B	~�咳�{�E�m���=̦��זG�������8�qHi�� ��0�Y���䬢��U6^�޻}���/}���e��!���e2�s%MY.b�8cp����Xj:cS׏5�n��9�b��S�^��V��������o�!+���5~Qn���wD�����6�|��2[^9� ����<s��������ř\���W�AM^	m</@S�8ͷ5��j�w� +�oj#K{y���m�����m�D@|I�L�@��>�@&��j���-�w�0w�]j�X��ۨ|sb$yw,����P/Kt)�k[�(-����.(9�g|WЦU��	��f��l�~͊y��7g3�����i$��s/c�\�H9g��
�W9)?�pй���,���V������UŇ�B%>�~R�r�Z(&.4mL��zr�U�q��\�5��t��l?v�]��<IߎC���O�\�~5�[~����?�]�ҷ7Po}R��V/P<��tiB`���,��A�t���[q��� �␋�?j/�Y���$_�l0"'H���YCY�ML<ߔ��c�7�"�}�y����*[
�OJ!�n](����콷����,\�-|�zxJ�K;�eB��2)�yӷB��:��{a�%�8���xl.�g5~\W�����6[�����܁�@M͝2����d�FH�&vH�������9�F��/�N0���~�, �����(�����ϳ��U���9dV1��B-1 ƳZ&8���A��B��y�_-mlD�f|�8*RȺ����Q3 *����sb��g�1:�g9K!�$f�kf�q��	�����t"����殧�6���8K[dҰX�p��M�0�����c�ܫhV(�J'�ܘ� ��y9+pb���B���}��r989M	IB^�~"ZlL�㌙vQ��(6�M%Hmh��jr��J���-Z��U�Ǻ�&v9�m��|��A�m�Zeod����#����y\��r��{O��q�I��Q�}�}���ᑰf*�'7�Z�d��m�j�̀�=F�7$��3fn��C,��T�|�y�C�
h�GY���l�h�_Qo04򣩹�&bc$agq�e��_�9*6��
l�U�-o�;��H,��l���Pg1p��A�V�*fBf�E{� 1S#�-��/f�O��˓3:�\ �Tb�a�	���G��U�M�gHfr�2P
����杼̊��8�k��*o:N�'��k���K9���X�6�PǴ��Lj��B[�N����
8����aĨ�(�n�ߨ>��DBf�֣W���K/j}�cM;I$�`�_�(Iy.8i2������c��S������k	�kѢoō����uuK��}�c�HT�-ȟ3�g�T<��iT�Ƅ�Z>�ǿ$�S���o9��m#���&����ԍ���ƱϹ��"�H��~j�����ς�7�P��0�2-ķ�䴎\�"�s�����*5\���q�.��mq��j	����.�{.�\���,8�/,�Z۲/0��f���5�\��CfVz]���=A��O96�~���W�7xͅ�d�擢)��Z��Xt|%�� ��GI 놻�i�f���xbP-J$�7��9mHhj~1�G��AS%8�h]���K���P�΃������G�Rbo���������$]h��+fE�3А�������	V/����8$�Zi����⏁�,�@x��.�$u��G@���J�r�i�b�Q[��V�������Vb����ɒC����gA�d�h�o�%Eeh�ue��N1	h��U���/�e�v����W���J�����w�w�Yۚ��)y ��>g?�P����4��؅0��\=�_��d�4T쯗�mp~W�J*����]�v����QR�g^�m�b|#e��ϕ)��3��P.f����Zj��.�ͨ�eh��8&���1HF����E����+u��e��GhL��g�q7�V둭e�竩�z����(y��1����i�NO/�� �B9�N��U�z׏��	P�T-��{|��ʎ0�q��$<��/%���՞Ţ�U��^�A�đЯ,����`9F��eV}�����E�8nt�< �Ac�Mh?<�Iý��CD �'(��R���K�@�����,O��|��
�Ƈ8Q9LF����(I���2d�/��!d�����r�2�����L���0| �$��k��c	6e���e��vm�|� �$S�>�4�$��%(��+P�eP�+��(���,=� +��~\Fm`W���~���k�p���(w�Ǫ[�ت�_%W�T9�^QZ�W�T���&+&/��e�A�
�v������_���a�-�ᑥ�h2�+�^d��Zl���I�Ur��q��!~X�N�]�0d0��|�Dc����lz� /lm�\�&1�ݩ�⢯��ТlϘ%|ck`�_�9���X�B�ƌ���SPt�X������@t5�~�P�^x?�5���$ȇV:j7�A�Я���Uֻ�_�8��g���_�J&@�σ��C�r��(����D+�o1m�]����p����mڬ(9�Q]ƒ���{S��'1�˗;[�7=�&N&�^\�(�D ��rQ��9�&�Y"#O���Q��,�R��b�d�J�O&�Q8dx�u��ڣe���d6Y%2�h���%f���+7�}�M�].��=�����8Xנ\/����6��+����=l�<�@ޖ'�]�
XZ	��A&�W�U��$6�����\�l�*��K�A�|M��ג�X���{vLO)�uҠ���p�_����P^���ր�P<x�����-2�&��Q�2	������t�w7D�jߣfr f��M�Ο��)�S-��.𔩜6]�qSP�葐_�!�l���5gVv ]�����\Z�lDphFUF?��s�(d�$�S��}S�� .]e�9!^�S��F�F���U�*�:��j�2�xl�T)S��;03O�L�t�0=��&����UG@>�"��sj
�*Ǖ!��)#�x����̭�طf��X���]�楮�{�F4�� ���.�zxvU&Jcї�1v�(_��!:.}��$��/)1dj�ǉ#�y����S+c��|�V���MmD&Z[fŋ���<$��I��a�]mc%�T1���cc�Qw"�B�*q?�f�!y�A.,/�nIGe� ���'͈�{#�:�v8����kr���|x|Nh�@
>	��Q��l`�5kUQѩ݃���6��Ѭ��-K�^�:I��}޼Z>𬷬��XB�f�ggfT�+L0SRS�m��q���&Scx
�VȜ/������`�:���8��an�2>�>�m�4s�z]́���8�R���(K�}a�j���u�E�~��d���Iӵ�m�v&�m�N�ضm۶m';�������>����ֵ�V��
�F�v`����5�g[u����־l��X�F.x�T`h�,Zu����w*N�Ej���� y�9��Az����"-�C���2�ܢ��P�9�h�-�e�����9��������'��c?��˰�[��a��σ!�4H���:�%�s��Dot��>�@�ܰ�����w��0��@��V]p���M�!�8�u|<aR�������^�|V�+� <�s(OuS	��� &ܸ��tyX�,��B�`	Vr�����޺ʋ�������.ؕ��P@�v��GK�U��P7�!���ԊPPY��n�����q���J�К��߲�(�׵��7���
}��.�3/�2��̦����68ܠ���̛	�X>N����q'���9�'�C��%|�F����_�v�od�N��V�˓�
����x����8�q/O�vg?��U?�At�G`~��'�Ϛ�/B��ϱ�c����֙��-�\��61��6#1IS��	���F)�Q<iq��W�2S�.2u�����R�
_ZB�֐��"�A�D��7�@��a��|����r����FG9J�%���9�d�K�< 臲������ф��∀�S���(l�H�2��1R��]�:���q�:��#�%���gq=-��\I+�7����
�:�)hd`�����xO ��vz�'UvҗGa�������g��������7p�|r��$-{yx�>�</ޤN5�\�f�;�<n����;�׌�\�!$x/բCo�EE˨�pt�	ԥ$&�4�ru6��j>㎠uGnu"�����^`nI�E��~1^�>�IGD�E�*	��u�r|�/����ɬ�a�0Z�@��Y�D2�]��Y�] ��rZ=�w��Eh��t�tuU|���*(���>�_�K��1�]��)�R!����{s�#�h/�uf!�F�g7BMw�6߼bG�~����7dR���՞pO<ű��`{nU��f�6՜Pd���o>�Oْ;��@�jC5c�O? ��$��Tl:z����oL�`�ԓ[�j�r!H��#�:5��Y~b
��Ї!s��R���������j*�xr�لPb�qj��-@JGT���"e;��:W_c��Y
����ե7��Qm���x��`�/'�2z�2o�k6"�d��نZr*����z��qCkyܹ��9a����CS�u�[�R��+��g7fr�8 �Qt��CE��(�)2�@|ЃaYhJzk�����>��|m	o@Y�O��qdl�%�j���S��.���+ �����kf�n�Y�N��f�e��;���&l��(q+�P��\��M���5X�P��QZstx,2'N#�xb2J�X���9S�rY�zft���b卫��F�q���&���b3z��<�w����\�E*��i6'�V�%�� ׍����؎ɭjgcF���~O{�3e#�\i*b���_[Q��(�M~�0t���}3���`@�[E��x���A��y�ߢ��U>��>�|�� AnA��.}%�\���h$
��^%��:�C��?D��Kvcso$�RH�UL>���P��Rݙ0��kCb���1�t�m��?j��8����0BIrP��V�s��e��t�A6�;��tMpd�>{	<V���͞�D�*�(�����%T6v�.���K(>7���?y�0X�������ł����*2z�>5+��`z�(_.���~���H���B�Ն����P���l���Dª@���4���&7�u2�Z�:�YG���ZZm���Z������F���/�$�N����4f^�BPx2Cq�9�R��`3�t���[ṯ1�T*aR�2���ۧ�~}���[��SR@� �VhZA�P��%��}k��}����Ѥn��Q�dn9����lo��1�������h�ȯ�x�j%�aA���J$�J�}_�������*Ʈ��ܶ5��<6G�*<*��/���ݾ*�*����א������#ƳG����roݑ�v�^�xPzH�l�1.�i�Rt�魆n6[0�o�Er�˓�I!��f�|(@�xb�����E���\�}�b��dR����{�m3���"k�TN���>����:��Y�/[`��_ၐ�.I��t�����Tu���L��������,q��ӕ�oN��SK�z���;��G��pQ��a?�""i4�h�L���P#U�[猧�q�{7QM�b������sA�]~��v�ڏ&�ũ4�/�<��}-�ԔI��J�o�r&.�ݔw����1lI�
h������x�_���B��w�.�q�FIޓ�o@�s���>��=:A�{�}A�\u9zK��#��j� ��{ϭN�٬.�h��o3��yА�=�B"8ix����v\w��ӹ�ŎD�d`}��A��.Q2D�y�I>��M<�O���,��h�
�cL��,��'�{Q2�%y�#t�U��FH�~!�Ai.3<Ϣ۝����<(%�p�(�=�L����L�q�����ɺ��1u�}�}�O���-�~a�0h��q�k��h+A��~�i��t:��0p5���E��7g %�.��[����K�n0L��J1�`��*>0���O��!�!�����19X��eN �����e���6��s �JF]D�<�<�"��6D�Ktƚ�ʴ%ky$�J�ړNn�P���\N�/�_�p�U��>�&�����ꌻ�S�HS��萌�V.\\�
�G�p9F9���9x���h�L���?O/LнG��-fb�#���2{��@�;C���Mx�VǑ�c��m�y��-�,�H�~���N�G�ݳ�7�RV���P�&u��|$�
Ey�����s=�5_��X�)�=����I}wָ���T�]{�(G˺Aʴ|���Un}_x�`� Vb>��5��'�4��E�#����b:��O�UU�:/m�O�hM�~�7��l��8|�c,�w��<~h�[0���Fgڄn3iݥ^�"<��hұ^7����i�g�,(����n>�o�_�	|a7� �l�@�#,�L�.o..\a�'��J�\[�����삯��o��j���r�$���w�$�4F ]�-�\��|��t\Ey��#�B#�%>���-�]t=hg���D��}D8U�=E���t��t2�r���~��n��m"�3X�N�W���Ў"\�ї8*Wx�3Z�E����%�^4��G��F3!h��wTc�Ⱦ�q�s{�un��	�����?���>����o~(M��V׼
K!`��	�����3k��/� ���.����Fy��/�.�>C�$6v�<��E���Œ�`=�ޏt�`������ղ��y���K��r(Q��jh/sصϬ7Y���u�uy�7�*[v�r�3�Kp[�A1-��!U��MR� ]�}���7�qG�q��ୢ��f�aB>�o_�=n�~��ͻQQ������:�eV�s�3@&�V{�|79�s�N+�m�>B���;������Y�ۢ$�4fh�`spb�WeeS�CKpz�ϫ_a���i�A�)�)�uV$-�(s��"�#���nN�6��|z��c��4�|t.�h�<��Xs�ЁĶ��]{��l`�>�-�\>�v�C{{D[~G�΍ �,֮Z���֙�~yq�������I\i 0>��I�,�~�n!���r��;����A��Jlل�����2A?��A����p��H�,�*L�d�AM�(�j�P�[湼�C��ß w8
;����0k�{TO�R|�矨� ��G�~�������FE���R@Ր�.�Y�\1���X�6����=pM�ɷ:�v�I���%��h���8$��[��7�[�"�q�΃Էt@�<ˮ���\B���]���Ρ�l�J�Z{�*e��K&�*(�tu�����ꠈ/�^�XеS7Z�g���K]��b0)�5
��q��۵oԩ[P���a�)�,��Ҹ��s�QJ�^o׫�P�>��9��t:A,����լMg�N�����ϰL�8�j��@e �K&�
C��#-M���1��"I�Jd���K�]������8v#2��	s�I�H*��t�ĥ�d��(�U�3
X�bm����Ǫf�A�ʀ�s�Ȅq��,��B��޸Z��Vc*S��M�Z� W�$e��,��qa������0F���V���S��g(�\��n��7O��*�.)�q�_���g�[&����DRP�d�m~���k������|6�S3D)~���L���
1jq���Y_���D��<����[�+J�s�k66������;���ۇ5$9m&[���KQ�ǳbvy�l�me�/���4�aÑ�W�Ԁ�ʝ�����/��{��d5��ƈ��!�HLS�}l�G`��O�E����rg/���3�4�S�ť�����N��͆�ݷ�mB��Jz�Cx�T��i�"Ǽ�r1��HT��أ����6z#�=w�L���Lp<��tZn��d����<��R���tC�}Nj+�^*�k5:/����#�T����,6J0V�U���������И�E9~�RV���uo�y���YD�l�I��X}���Y@�h��r�;<B�����^�N���ÄS<�Z")�Cr7�hsH	�m&) �8����ƴ��YpӷbsW����԰a�υ�Q͜L9HU�PN�dR� ��}i�dZUHݲ�Z�H��ҭxxQ\�10|��zD��7�<��C�j��xn�{���E�m���'��L�i�m�ͮ
���Xq ��T�r})��a�>��N��nO��J��8RMd��t��P."��3�C]!���Q\-*�0�?���Cbn� �Mc��K���稂��� ��|�N����1��(|�o���t�+�dE�(w��r���y���*y�<�[��5�&����MW�AIr]}#����0����2�X�Z���������Q�le1�K}���V��`8�8��r`�n|d���:��Xc6��e���weO��_M�Y%����Ƅ�����V � ����c@�Q��<<C���l���*k��� ��̐Lڑ� 4�(݄�!�~���n�����9��ŚW���wg�@Ic{>�:�:F���b���O>� �;W�v�S9#iWl���^�T5�#��cC3~�@T����ͨ��:&b.?+]��Z��W��(+��z8�T�`ϚuK��	M��C��4̩;��ý[�!��R�����ⓞ�e��e����ʀR����%$Y 
�i�Q�)>��Y}t`���w���dU���Ms�d*�`��2�)��:�B7�
��QI�ң{�m�T�dh�uTB0�J� ]�'��+<�$�Z��{��;��G�Kc�yf��L˷��,��|t T�	��.����JI�W�y��zQ��7�7m�?3�	z�r��	g�?{�ؙ���x.&��Qp�����o\��N��������U��>�{�0����A;'!A<��;�o�D�.��4������icq�Qp:B[l�������9��T�����Əl�a����,R��o�Mi�3<��b}7���Mz�&n�#3`�Yl���[ә����"��i;t*�,��X�MO3Y욢H���k6�I��X��ո�F�\����0\���K׹4�v�ibB��B~�@�AMȤ3*2��42 ������(��G��O*�lve���}瀖>����\pP�F�bo�ORcW�#�y�K �!_T%�?��r����e"j����-k���S�إ\-���|���S����U7������s�op]�ɍ�h��`�2��3�_���De�h���e/BM}�卟W�/��D���d���[:-;�Ƞ�K��f��Y�����[`S�ePu�l
E#�}��a�ݯv��Rf��ph p2���E���*g�"��J@��x4��K�g"Ai��+���-h�48�1fft�b�Y����OuQ`h�R,�.�}W)`7�{��v��Z7L�{�b&6���Ꭹ[61��Gm/�]\�Zr$d�<�Hx�lͶ�ͪ\y�4�0�6FG\q����8l�fj�����s��>*��KB� �{e3��S'�4�L��a�eD0_��-���w�*P�8��'�l�Xv%i�(l�9����n�_`�y�͙��<{I�qȝ��:2_��W*1�o]�_����r�Q��#r��' �qN����i󰄶�"�ߥqMb;�����M��l\�T)X��@@�$+���,������ڼڔYifʯ�OLr�#���haZ�lvW�t9�7q����@�G����e��^&X1dv�))6 �<�(K��8���a(�>�4p��w"^=�*��k��b
oM>[k�݀��m���?|��F�*�n�VmY�46�+�gf/o�f��Ny_�+��Q��4H�l��jZ�X� �k��a�/n���-5�Q�#	��I�<D���2[�=x���~ʠ���2�����lm���sǵGƀ��O���p�ɘ�-�)b�F�& ���3/]��JY������x	@W;d�J��:
Q���Q��tM*p�ZόS�Z������8 �u�m�����w��A���4 a���W(� d���5�<t�O�V{K��ʑ�C�6�}]�3��cW���vc�S��CS,$������Ud�I�L!�D��Y�m�247[��s�!��틏B*�??�[X	1*irB���PK�:����d�y�B�q|5'��M�OP��Sg���~��'#���cL㌗hs��8�Goz��G����/��=?��G��x p�q���C�W�����`fY�!v�"~��[���<<+c�%^ԓ����;�*�5n�}_O.&7	���֛\n�}��_��e/t]
���>�4¥C/�Nݘ�^�f��x�v��"�o �}�>1Dq������{�������jԽ�
ٕ�G�o�K=m��w:}��m���-�M�aK����O�մm���s�NXRK�|Aw�?�|((�y��ڕYLupܤURa:��jߴ�y��:<	����WW���E��y�1n��ڄ�i>i�(�G��xa[�.&��&��QO?��T���>�e$�i�7�� Y�F��=_3(�0�h_���-�����&Ҡ�����P�,�N�L��N�]����.a@Pr��hN�)d�
9��3�$��%5~���O�g��Q�3^䋷'�Ћ�K�I�%D��]H�LO}�ʭ5m���c�,��|O��C-�o�e�"�[I��h�A����+?r=�4e�ߕWC��g_>��Z�+��k����v���6͓uK'�c�Ww�N�:�I�KgO��۫�ck☙TD?�F�֌��;�PH�9���^�E����^�Y�Zwz :�0�K���V����E����:H��eZ�{8����Gm3�H�!r[��4~����֭�c�.մ)�\���]�y��������JDD�g����ŵE�z��r���`��~�(�|$mF�ªQ����T���/��E�I���GvzGR+�E:a��T�J�I�^w��ºl:�G2������DQ�K�M-�Yhn����wۥ��e/31[8ENR�А�T�>��?�nҕ�W#�߶6q��,I'��'�T	�M爔��U�ȩ�>��Z�?Md�܊]�H������y"�Y��UCؕ�Y��%�Q��&d���bE�-�K��:���\Аdv��������Ndy.ռϦ� ��IgDJ���+U�ˁ����ej����CO⫵�f�T¦K<��BEj%�P��As)ui>�u�
a�Q� ��o�(ʻ)̬$AlE��)����Gu�I�]<�0u4����H�&IU@�'�9�7��y��	
wQA���P^<��`���zr��R�%`�r�����������\�_w�#�;z$4�=�T���U��Gf����E(AC& �8�A������py�3&b	|��z䙘\p�"ަ���Lf ��a�������b�;�)���T�u��L.�ѕ���@E>�O�LV�CSJz�	U"moC�.������zR��ҙ@]%��g0�����+�ؙ�IS/YzɋRA���ҝB>r}fX��(�~o��{y��YFn�in!!�ڰ$`�4u���L�-
hB�
L�Ej���nA�_�Y��0�Lvc�ι����H��׾
J�����%x}Xެ'2ۋn��F��9J� ��
�}��{>����O�p�Yj몒�\�E��)�Z]ؾ�:���s�+��}K��M�BԹ�U�[i�q�@���y�8���\�"���9��O�l�zzChF����X�xqFq��mv�`��M��Wx�I�Q`���;w)�^��?�דɖP��J�w��L=�;
 v:�6��ϟL��!E��;Dl ��Ĺ0�ʥ����3�d�j�nD��Gl~)�6�S�5�*8熻)��n�f)�q���%�R[���8����5��L]U%I����G��bԥ�J�c�Q�u�M
Z���XAi%hUs7��������x��=�t)��������D��?�-���(+G3��_6�5��������S����fx����3�����}�_���p�~�u�����gIn;Q��� 0E.`о�4�	Iݕ�9q�����C��iti�5#?�Ҟf�@���*Z٫F.��� B(��. B5Qo���y��dV��"�Z�X!��-+ݐL%��,�Fo�ݠ�J�L��.�	ϯw�C̠,͎�,��Iy�U�L��{�./c��^��)%-��I�.�4'�h��.����	�dR��hn��ŚT�#��V��!ۧ�(P�V���0�?�Xz	c�_0�(��x2łl�$��5լ��m4U�SN �v��ɲ��ɫ��|�vH`�9S����'�p/���ua�c�sV�jP(K%�j��fe��-���4�G��#΃l��3�u^�>�m��V%��n:8޷P3[�
��͕i�Rǽ��f�:�HN������Q+��F5Z�ⷾ>1�ӲK1c��}q�tI�*�2��a�Ź����C[�~�d�`�o�oX�݊O?+�����Pl��2B'%c�{5u�)���BC~��0gv;�葕�_�l	_�K����8�0ٓ��4�-*���d��?`�3�`S���X�T@�t�0�tc�Q��$\#&�0iޜ&�(_����j6F���{!���5���k	'���c
*��I�bB�������1�1����+!�iA�pP4Ϫ��gZ�B��XIs�|����4�w�֑+�kߙ�V��@�ǫՔ�<FV;姣�Н��z'�dE�UԨ�y�����*�O���M���RG4�{)L�Z��J�[�I�AbZ4�����V�3���ۻl|�S+־e�1��1����N"H(���狋�UV��~PRS�EϳQ{\Z<_z��9OWyA�&Iդ�}����?n���~A_�3�E3jat>�~3�6|���#o����=�D$tp.)˷�w!��g� �)!o�1�!�/;�G���c���ʴ8Q��x�1�bD�������P7t[-&"P�U5�f��B��a�<�������)S5�!G<����#����`u��뾿J z2a�
��k�pA�����������|X�R�dE�b���I�2"���N�-�udsdnaRӢ~S��� QR�
��d�����U򣎂�������{{����>dƞ2��͋��ۡ��hA}���USk$N����Y�{�`����p2k0˸lB�Ms������~���^腊�~ϒ�PKɆ�n���h=�!e�.�p�X~}XA�$�hac3≼���Y�~ 1i��`�^���u��Xq������öU&�������A��J����!$8|'9����D�5ckk҆�.����)<�F�iTh�gvT�@�����g�+�@u���	���U\e%5�^'��8yu���n��K7y�ղy��D]mٛr7DT���S�{���y��0��!S��5$7n黉�5�6�j�86�v���nT�9�H_����u&�t�u���+�+�k`K�̈p��������'2m���_3U������������h	&U��̄�zR�EQ0::ۈvOE�5�%���F����[�U2�ݢ�x#�(�g����cc���3 ���*אB]/�!EM�3*ר�k]�q����KJX���!~���;0 UVx������77�v�a:�A���D5�YV��R�JH��qwޯ!=^��祘I���It��������_�� ����3���<)�_/[��j���i0.-�d�X�G@b�s~�ꏝx?��Ef��YrO��5
���B��r�X�.}�4SWtN|����T�@w��b�Ց%�`@b_��o�GEE5��t�ݛL����[�\��*������l���y�Tʷd�%i'�X�̞��8����vt�)�x&RB�yGHܠ�uSZ�ζ��n�$"Ur��Ċ��l���@�ӑ꺙%��T
7�7k�V#r��]n�8���IV��^EҤ��U��TlkHhX�X7R~,��'<�T�~�b&�F!��'�Y����#ʙ ���̻!s�oډ�RRQ'�D��"IHwz8�#Db'���h��̃��t.}6-�.�}@�	�1��WP�E����<21?(B�'��$5�.��bobn0����:7N���S�d���)� ��S]SU���O���+�H�����u~���ȃ���V�l��h2��l}�AN�cK�GƇ�v�iw@����L���O�?驤�.�����4aY�AB\�r=>V�ZgV�֍`�V+�����}�# �kut^ꔷ��l��/涒��<f	���.D4�bQO9�{,��`�'��ӥhˊXw(���H7t��V�j]x�I���zEx���@s�R�_j���Kooo�p�����(��V#���8��5�B}�z?�a`�8(����:)�g�6[�@H@�4:Kҍ���0WW&�;��w�읝��~���!��?�t� xK���Z\.V������]?�A�6Z(
�
�J�g�U�����{_�'���B���x��**�ĉ��wvv8����F��;+�L���-Il�k�f�=4Z�𺿀�R�灋�s�7�y���~�6ۆR ��rPX葥�3��~�>2�|��g�߿�e�]>�����J�s#N��������@h��;k�\<���z�=8+<���^��|"��8䢦@�_\��N�}]cl4G�b��,D��;jf>���,4��/a�@n�th'���4�����U.�
�l�Kt��0Iİ�4�"��E�=?$ZP2(����Ԇ�%:����EW���

sl*(�Ŭ�u�/+��5D1NvGG�N�Q����STvG,N�#��)��$�n�?~sz>+�WQыi9V�۹}�Ț��R @�Kf<"B�IEx�H���]9\�2#�^`�?ZS.n�Il�XG�@���Cj�XM��i�����|ģ�n�VTT�_,�LB�].��������/!@B�} ��"G<;t�NuD��Zv"�"�Fui  �z�<�jГ��I��~akGv���������qI��@J�����
w'�O0^��E��F�qCp��p�JI9b��[XJ���c�%9�b��z���TrU������PI��}��贎�dG������X�8a��) �==	�rAuC�b}IM�@j��bi��0�S��|`b"�5�c� A����	�h]i���K!�Q��?�1X\V u2�YJJClaf�����wʘC� ����tL��BAA����KH�m����G$;�һ�� ���D'2nH�7��v�4�]Q3x�7S9I�gб
�D�$�v�l�|���[~\d0H��?QD|�Z[7O�_��55 ��SN���d-�t����J`�R�	&JZ1#�0�1,���ery��j&>�[��CP�
��d�5�s9���Gd:`鄫����������Fη���VS������h_GL|��wB>Litt3�i��vŃ3Ut1a1��)�)�$�~M̶����	�K�����VTv�!5������9�3�2����Lm)�2��G��5%�Z�=q�I��&�Ԟ���۝��]�\c��1��xI��m�o-�u���,b%�p�M��8R�U��������-˸>��ax�����E5��_g�.�}%}�ݚ���.%}��>��6��B�a�������T�}v�5P�Ex����(�����R�~���{��@<�D�K�տ_0J"�Tk�����)��=#�������>�3��K��4x��I3L��`lH�v������aYƚJ��Ka"j���w�����w�ZC�U��ou>ܙ	ʡS���603&��ydU�|Hfh�ݬK�������two*
K[�-��\{�-#!H��Lw&iL���j�oOj2m?@���)��n�rY��i�:���_;���ʺ�=�߂砾�ih����J]�p��.�����en�5eR4�I���*�MJ*���ܰ�ޤ
X7�M��v���i��#V"�:b���[.��W7\gv����2��M�>]Oe$u�v:^�N��n��!�t���n�X� q��fI:�s��W�����4�����-QF�*�h)�d�t�I����2"���[`���� <�9�4���8��{^�]�Gl|Ph|E�FiVP�sbB��>���������~O����s�q��F�/vt
T���}�N�����������>X�ؿ	Gq��w�j��n��K�r��c�W�3��@�~�'>n1����R�Ǿ��c�A��-��;�|�G��@9���#��?@"⇀�����'���h�d�Ҧ�3���J�5e��1�c>eE6���[��g�e�+\|�[>*E�b����GO+/��d&(3�
� �������^GV>�'��|.�c�ǚ8�Kq�T��q�X���v�m����#����k��y�������3x6��X^����Ah%=����|������)R{G�|`.w�-��r��D���4c��C��Ȃw-��U�9#�Mr�@��u�b[&�7ȩe���5E��PRc�rh�3v��GIM/���?1�˪�²:�(�$>.�q�y�ʥFk(�h�
��0�����I�&����̴����J�P�����=�.�<��R685B+n�ތ��2�y�v�]��� 2�VV�� �G���x���� "/�A�F;���(
�-~�����������-���>E���fZ�}!�������2L1��5��#���\�.���������
�T&�Wf����X{�O��I�,�'� �r3HR�,i�'<
�q�B�j��rnqS�f�݊N.'��5fu�O�qt
eo�Q��n8I�	)b ��敂bpDW5�/47�y���i9��q���ғ���]d�{;X�������)��v��v\\f�2:�U�����NQB|��B�Z�D)1I���_\߻�hz�ީ���=� �Ԙ'py�����@_�S�����yc���ix�b�=Kӧ��{��Y��n�ho��_����T��K��R�EL9�YJ����+�R~^��[H���kq� �k8�Gܼ�͂"��?w,�
ߛR�=8��F�81��աB�dNLO�.��#i�)�@06�M���/1��>5��G�,�B��F;��/#�<b����־�J|�ߡ�4�n��Y�0��u^?Y�����5C���t��oМ�p�+�����G�����A[���<��L���0��v��'}��2FC��!�դs:��6Έ��t�����K�0^X44"��x�I�R�������5�T�
?�>"�$J.���<���ބx|�_�Yb�,q�-�jN��?,L���*��\_ĭ;��Ѩ���Z������#�:��f�6�_��1ڜ*8CC��u�R�����>w��x�-�oȆ��BBE���P|7�Cʸ�Ic�*c�)�d1�Xt����1�y������8�����ԥ
�A֞�V��	����>��:`?7�싖�542d���U$�n��&q�(�e����T,g�i�G�4�?=�)�K}�[b�։���IEJKb1P��8mO˄�Q�1��47.(%����Q�_e�&���}�( ����$P��GFE��p����D?:�Z-��������F�����D]q� '�i����<QS�`Q�MNJ��[m�H+|�6�02���p����%&X�$.����F��;5{���̏�5^b��lN�-k���eQ�_��R�SL.���'�
�jk~�^��^Z�IVU#�(�Z�u� ���.�E>L�Y��Fp��u�/DO9:���� �����IJ���w�&����pm�K��zF�L�ppמ����i���G�����ju5|a��,�0-�򜚉����R���г��kg�����mbS�WW�y�L�&JjX����@������Ԯ��]��.�ҽ�:q4�D�l��Ǖ�V�km?Q�����%�}G� 1v����rQ�2���n[���*���f�n`��V>��;Wm�)�I����^!UU���ឩ���4���&����V:G�]rM멌�4�u��TO���Y�1TN�]-:�</nq���n��M1�b�!`��ź���t�<+h����mA)2�l�Zʓ+g��nɇ�IH���3�D�7a�Y�����h4�������r�Ė�L��g$�E�����\����^�*��Lm��i�Q�I�z��/9�HZ�?����g;ք9;��c�O=V��g�ί]�v�
̮�����a�k@��<~�e&���w��H�T��vz�����ڶ�|�L��i
?����@�t�n�gDl����֌����O���|�AW�g9e��N���T.��T�E9��O2Vhhe�Z��������%ϯ[O����L!y+*��BY�{�@R�f��T�����-Mc'ҩ���ॣ�*�F���H�դ��n/r�������>Y�QGm��<�}.�a��cC����6����	�b���Ѯ�t]���c�q�L�0��B%��^|#��x�H��E{����;����W�~W�dr��n7����^�A^�f�9Cͩl=`�Uli���Ӂu�⢂\�B���$vpsU�OUu�` h��]^6Z��O�z�N�஼�y3�َ�43�P�����J��qN�|�+~�T���a��:¾K;R�p0/�3��B�ڟ-q9�T�y)Є�n���G^Ѝ�v:����6�(A����r�j�����P�o.�7���w���ٰ)���𨒔�tb�[�S��lW�aN��?���
&i�x=-ɔjT�B�<<;>��j�6����S�}�H�f��<���AD�ym�?�-P��I�D?�3$���_��r��b�l���X��Q<,����E�uwwW^[C�h$׸ABL��%�V����r�
�w<��GG�_a���$|�^;�^�|#�Y��NV���s�v�l��J�dE�Z�	ʢ+">�>���^�ץ6��̤��R�1�&��t��OwINL��j�������T�3P��I�0�^�>����e��g庑�.�wJ���r����=���f��H$~���Pfu?���(��=-bX{]�H��X	��H���;Ǆ �pp��Q���wR��������q�븶�A��)jb��PA�j�N�������u�O[��#-���+��kB�.(,�w���=�KK�Wz��N	�'�~�p�ŌR!u��
Wai���$�o]�,k]�#v�0Ì������,��x8�Ҋ��R���>��h���'�(�M���=���C��d�p���M��_YW̠P�`�s���istd�u]����b��5;�W��S��~�<��A0�]�"|���
z��?�[E	�Lw�Ʈ�Ӑ�\ޝY-�a	8�����J"�k��e���?����c�n�~�`N�WwX�F�i$�ߖ�l/��1�Ρ�`}v���)�7�m�b���d7D���X��1N�����p�3�1�_�03-�~h1��`l֛L����2ޙL���`4o|���g��_-g��aN�CP�z� |@��
�0/��������C��c�y3KX"y�XiIc�����S�bڢτu�"�/�������0�x�P�T>>f�8m{��I��Ԥ�ѽw?�����٘����L�zR�_���ָ���A+b=|���ٸF�=rӞ~�H�Ƥ�s�����x���g�S�f<�6�:jʅ���D8�aR�r�'j�<1^M�D�������h�F���՚�?R�'�d���{�ZP|��%,6QQ��ҫ��c�f��/�f�X|��"��?���v��xV�/i�׭',�M��'��������h1��̙�뤱���^��?|O2O���M�6UM�>Dl_�9��+s1~�x�]��k|L�{+�÷S�8_|��~~����0q�d�#���:�94m�DL�6C��\MraW���V�����1;��v��[1�G�V�1!�N����Ə��F�};o,x�=j����p.n^�M�[�����q�����h��A����z����/�W^À{�#�{w������t멩ϖ�5��o�w�D��w��T�
�w�������O���侢s������ak-��.����MM�Z�+b��:)�O�H�� O_?�gܠ�q���#ZնV�.�H�����ȿ]���r-ҦB7O��rg�o��7�^=���3,,,�OʑO ZXZ�R��k뉚�z��ڗ�N� E����;w�A[R����}3��vo���g�B��.@^N�iS�#}�w�8���k~>ro�CG�����(�9�T[ww�?�E���h�V	wa�`t	�]�Ȳ_@�p�wso���l466isjQ_۶�053C�&os��ϫ]����x���Q]�@m�n��]�bO�nqZ˗�~��y�ղ��`dhJ�uq�x���M�� ���L<�\M��C�v<n�s���E�bd���m7/__4���C�Y[��u�?T9%�t튺���n/���e�6��w;Q�εo�11g�o�ڧg��>akm��p6O���ë=�--aeg#��j�o#B����w �Y[�½���.��g]���ϥmA��ml�L��)��۷C�r�nnptt�����]��}Ӛ��yX;8�����;�D��mn��qؿw/�in��lC�O��r�++K88:Q�PR^�������K���gE[j���ɲ]�r�v.�@/���Eyy5�]��xn��O���z,����?^��@_���o���Z2���
:������ј?�Ӓ"��_�0h�퍇G>VX�ԫ+��A,=<�0��D`ԀN�����j}�۷Ô)S���H�۵Z.(�na��}i5��ߩ�r��Ï?�C�^�2i��+,ݮD�ؚeE�)8$D(���J��������Xq�uǁ{O+kX;:@�ФE9V�.�L����\�p]/"�O�W�EJ�OC*X������+��������hg
��C�?'7��X��v�:ء���-��cKt��o͛�j�l�pL�6>$���J����1��7�zK\���믾�j}���2j��*�h�ÏjY� �������A��$e�d�lmq���s����-���&hYq� ���s��� 2)̞=W렍Z.D���)��(����)�f��5F>�y?�`�K/K�m����1y�R}ܾ��gY5���¨>_"9�ֶb�Zضr��fΞM�ao�L�Ҫ[[�{�qq����fӽي�	3�y���h�o�{�h,R�C���>t�E���#H�[��g�G`� A��z{�D�����=��^b.>1v�pUh��|.D���O>\H��g�2,�aa�$"ϧ��=o��h�(��ϭ����
�uC�M	�U��ߊ�C�2�N[�����z�w
��+V�Fy��_���5����=����~m��եI��䀟L���Ш�#��Rn��s�����	 ��R}ϟi�7��y�y�����$����x���-T.�"^�����B{�j},9ն
�i��Z�!)��>R93kkxZ�J��=D2��Sj��=|���*�=�K>BL�Z/G�3�Go�'�Ѓ�&�]����#bbe׺���T�N涎�C9�ʒ�JOsJ���3V��c�p��Q}=��0V�a�^)`�&ޓ����NP�N1��m�٠��rv����_a9�m�֡�N�(p��������ίk�
�������X��b�/��˩�3&�����S�AH��w,��E���~S�_��j>3�RlA6���!��\.���Z���c9e�:�y<x�W�.!��XN9;⯂��J��aA�;�p)��dh ����pc�|�뵪�T:��3�r��;����&~Mw���қMw�պ8n�p���T�^���P蠃:��׀�U�h�b��S��V�FN��%}T'�W���]����Vt�����Q�KF:
�n��e��)���/,m:蠃:��`�V�� R�DG���i��Q��7�5��88�?&mНZ�At����6�F:��O�*��
zr�G�����O����(�j��E��At�+�/��������7C�CO�H4���N��p J�V�:蠃)8.��<����ӊ�b���o
��{m}�%��o�_�-:�(�w�Dv�M��gȐ��۷��s�����͛P^^KK��vĤ�Sa�,vXt���
GQ~��uxwϻ1���`�ߌ�@E>�\2K}���Ӧ��q*�(��م��L�8|���1r�ðhD�\�	�[��E014�� &L�7�f������e���'N���v�ۓQ�����`ieOOO���۷Y}DV���[��k��x�������@<�ׯ�Q9s�����G?ޢ�c�U���DUu5;`Ҥip���z��A�?�_-���#����J$&�cŊ�QZ\���Zt
��ɓ��,�V��8��\�*�

�Ï>
� ��z�g���Q__/���u�iӟ���g������i|sQ�P�����8�����<$'&`��(((s���*:v��i������'��� ^^�;~�O;<G���_��So���]躏�z��uΝ�����z������	�&�oQ.#5?���RSEN�v��a��a��S;��Ջ	ؽk���8|D{o/<1~|���HM���kq++[�krrr��M"���[6##3��F033œON�&�������#����E�m�1��ܽYx��t�^,U�Ss�W��v��Ӱq�z�Ĝ��upĐaCѳ� �r�9YX��7��9_��D:�G�������-ԏ�i7PSUE���F�����fga�O�������F�Z[c��0���V9�� �J"�
�ю��8{A����#�74h5������L\���,\J
����<4�������ܴ���ůY�~i{�N�����=�Tc��է~�B��;�pk����<�MR�FMR�?��wb�ڵ"����xhœ�_���{g�����0�8i2�--E��S��W�B���r1�#�����������A����SK��o/�H].��C�@��`kq":k\�g_|E]��'�Q:}�4�m��*ğ?��?Z��?�L]�$����}���&<H�s���q�X��G�}�mu9&E濋9/�w��ⳳgc�����oi��~��$��ptv��O�8��>�K�]�.�_~�9&<��H��qҸ���W�W_���D:��m ��s�s��x筷����Z�-��c<������ںz�l�w����P-�܂�?��ٳ�=�GdW8�<�{��ٴ*k��EL�n$ڷ�99Y!��Rj߫"�#=�*^u.f͝����`�o��4n/���U�W&E���2fΜ)r�VUU���濇O�,V����+xi�,���"c�����l�'X�j-=]����������)Sac$_��e_/���>V�/;=oP{�L��A�	���^ǻ��׬�gD&�Ξ��Tߣ�<&�N޺u˗-���O�)�`nV>xg��<D�Ђ�||��C|�t)�xu�9/<O�sF�~T��|�"��+|�n_NF��M<�P�B��D��ƻ4�-Rg����ĜY�H�#��"J?'���W�n�F�҉Q���E-�С�1b�я��\|�٧��O���T�՗�b�c�02�a�ʊ�>�˾�U/����?��D�gΚI��
�����g�E@� 9�^me��1]��z䑇�s-��"�+h�����773�����=*(gIټa\�]4i�k��0f�X<8�A���F�qݺ���i�θQ��+�Z�n�x��	�|�����m���� ��xgޛ�w���4yLMMq33�W����-��A]M��w�}��m��3^���聵��X&�Yϵ&s�����eq��:����탷ߞ?�Ղ�(qBt%�����߀�"��o_�{�-��C\e�wp��%��[�gҁV�ӧM�Dq����,X@
C��g�	���8�It,$声���uǌ~L(UD|O/O�'������-����j�'����W�"Hi`�pOL�:M�8�����{�!D���r;�62�'��5}��˯hh� �����>�Y�:��mq�;�~�n����q��."-)Q��]]D�IUq[X�w��Ϩ[K~��V�||;��8�����cҤ�D�T8��"��-��������|�e���C��4�&��'��\Hr�\���C�F�TV#GGQ�r<80lj�5�=���ݽ-> Bڥ[u9���E�5=d+���^���B�)8��%�ũ�ell��罣5���gq=�����u���/`@���Ǣ��F�Bd���섧i�S��^�~\!"�OSssZ4��p+���s_TD���/Q�3@��e�$4��%��/]�QO>5�E�ݟ����ׯ��362�s����/�{�D$�ϫ�w:���`�|�W.%���R�7�~z�����3o���&']U�{��n<d��=�]����lq#�?e�T���\]���34v#��lmm������$�B��������w�`M��p��{3��_B�t�w�W����n��}�x�@G��Qǝ�|��b�Rm1R1�`��'�4rm�mŰw�#cL�U���j�>#ZIգ��HM�:���oe�Z�W�U������x)ad` Ƽ��ruZ�SCc�zk�׬�9/*���ke%�����00�GK[HO�����)�Tpt���051E~^���y���y2 c�窬�մ��Q����Ed�#«�D�tjv]+c#C���b9F��|��5�Qh��U�MQSS�����]�Zԗ�����:��9���uu5�yn4'mR9s-�p}ZIJ�sP_a��tWJҦ�%���B��l�vl��ÊvEY��o}�OI�T075CY��[�Z믋�4�}-�A󠶶u�r<��%a���BAA��}-�����[��
[�6Fɸ��B���lm`e�I/���J}v�0*+-��LI�Tp��GYY)t�A���죕v#�܆�xH}�J��1���(�=+kK>f&f"	'�V����L#%m�a��\�ZC�̌5�y466F��q���"3��r�ݿiii���F��3�<�ǩ��!Æ���V6V0����۾�i�	ȇQ}.^"YvS���'���g�F�o�a�`�Zkg����ˉ��"׻O���-!���Z�b�#p.��؆�{Ot�,��x�Y�s��q��)ខ��tA���Yj�3�#q&&u�ub��' %��85�V}1'p��q������CX��c؇�J�E�Oj_�.���9N������u˫*��v����ئS���###QO$�A�W�֊�w[Xh��r>)�ؿ� a�㼩�]INFۨ�=��@�
�	�q�|�ɗ�!\)�"�V������Ç
B��{��Έƭ�T� \�����hq�s���;h�;=�4���sgp��Y�R�BB��"o�j�Ť$& ��a��עK��8t�xc��k��^�z?o�
7�P�7>�/.�no7ǝ������r����+�q=G"�£w�����i�fyW�����C�Z�ה���;�������ǢPTT,�}/���5��/|J92����6#Z�-}���Q?:�r�u����&�9�C�Gyy���Lp94DI�6��Έ?L��N�x~�/Z�Z{H�^D܇;��m�;w�S`'xyz	�n(1+֯͟��C����ht�����������
L�v�
'E�5k~D@@'���%ڪTtLb����#�ӆ������b�jW���?�Ƹq����ع\۴�����ڄ�Q���/��}��hܾ}^�Y���Q�����'<�uk� �KA�
�h�hny&�K��
a�D\�yR�P}��Ny������/ǔ)ӄ#9oM2qc�DM��B�����Y��g�n���A��B����VC|/����K��C$����Û�c��VH=E����S�~ٷ:l8����G�3���(�tʕ�X��3�?���k)I���k�����%�4iv�����	�'�]R�:)W��}�ƌ��#�t� nv�v���֔KM�k����_}1�N#))�D�jQ_�!�L�>_��Əǉ�HINĭ�V�D���G.Ĵ�3��g�{z
�OD�N'#�*^�;O�xǈ4��[
�VG���͟�"By��5��� o�s��}�9�x��y��DB����"ä���D��G����)�f����kY�*����o`���HNJ��/JiY9��u���<|��g:|(.]�(B�0!�1��0��WZ��O��("�r��^5�SZ�؇�o���|���[yik��F���PX._�������ZYZ�J��ZQ�������^�D�c��3qc��P���^�;���-�9��_ ���d�b<�ʊ���Ǆ�u�31�\Eeթ��|�q/(�~p��Q}:[�����h;����?R"w�瑚���#F`�0�<"���YX�i�2�I���=��22ah`�z�����X��/i���a�"����u);;;���i����A�Ä+..�98�iYd.��z���Bj==�p�6��[�R�(0��	
�7���<��%⡼��u�S}#������1,,̵,x\G�^�1j�D��΅���h?o�5*���T:Tl��:yLm��-AS�VЍi��zaə�},�F�P�A���t"�]���|H䙭m嚭�|t���c�&�+��lz0"2��T��W�@%�ݼ�{;�j��WZ6��;4��خbYZ[��G
��$d�7`kg��QO2�$�b�ç�娿��۴q�����*q�|�=�J"�uu�2�f33��&%&b��{i�ƈ��ؠ)��/';�H�=��M�Ҕ�rK|��2�s��/ ����U˾FY�f{�O\�PYV!�"G�� ''�={V|^US�u�;7;m���x<�׊S�GG7��pjj*ڶ�ʱ�6!��ܔ��~�*d����m����2+���@�
3+�m�"l�8Di�>vL���B5w����̂O���4�$-�,�)��ZXZ��ur�Y�*+I~��

�r-�~Jr6&�$���\�\���E���ѣ�z%Q�`�i��"u�gc����"�8-L��c������}�N�F,FF=�[+m���M�.��GN�������M7N�V��8��g�wC#c�*gb�o"m��D����B��[X��RYy	�d�oV��Ũ"�gBu5�R�,-C�,%�hF��::���%��F����P]^�n_iA!�H�0�*`n,����5��WI�H�l���Ņ�d/�����ϻ�C$L��y�D�[2x�L��M���׫�eN�U����Z1lH�W��L��%���r�G;�I�(-G'ga�`�����*��"��l�8?5�̆�ZX(�QME�l�,���.��bl���+[J�e\)�*I	�����]V��
V���<5*|�x�eRr;7��KN�lI32�(l���L���`/o/��¯��AS�U�X#�9�
S_U�
�ϗ��%- $�P�m'9�A?�5-#Ƕ�N򵊄<��BOay�����L\���<%��Ra�Ҧ�N����F�ol��+�i%����2)��Sok�e��VC�ؿ��M���s��66��Ԕ3�ׇ��4k*��h+�&Կ�j�E������d[Bd��RZ,4�Xh䒛s��K�W��]Q*�ր`J7[%��\�XS��D��65�5MD��Ȉ�"����TS/˲��@s�UPۍT>rU�ɹ-�������ߒ�����j��ffR�)�D ]\ڠ��G5-�����X)/����Έ_%n�x/:��!���g5�qqmC����Py�pX��J~��Ú[�ꈐ��p�&�J���D�<���� M��&�������g�-���,m��Z	�bl���1�4�����I�WVU
�h��RnmVу�^~��v���}o ,2Պ�Ckk�0��U��	[��N�瓅55�|zA(�[t��$E�
���6�6�M?�Ҕ��*�yk�-��,��k,<lM)�	�I>�+dTW#��7	122���Tq3S��ʂ�Lи>CY�������C%gv*�o@2����}�T�S��9:j�۫V�z&������N(m[�L[�4��[��cE���UT��-\��nd$���Ȕ�WV�2yV���T�j��5�6
[۔>�l�*��e-Gk���%���*�e�\����m#�2���D,4���c+tJr�|�0˨RȒ�dgeIץE�������b��*�:HL4���[��~М06���T^�����$1���\Z�����	��o��`�!d���R�R�Z�0��QR��.˲J�g��ġu+4�ׄ��*T����GiQco��g<�
�^�CI�u�XP=k�Z�������&p�R�HMUh"����Yv�P���uk���GlձnT�;�t���i��k�/˷��,�?�ïĉ�A��=�c }���I����^���N�՗v�c���ZP^�m)旞P�u�Ł> �4�~�7 ��E�g���L�1��mLzh�Nl2�z�ǖM�`k��qQ]ׄ˗����7);��rG�.�i�z����KK�k�\O��v|y�P]Δ����u#n�r;}��^���=��a=�"<|'=��PF��X�Q$�$����.�e���qd�Z��w�U�z=$#_���r����K��{Qi!��ف����?h )AM?��xcپ}h�uN�;�k72p�v
J��޾����g�_�f� ������oe!(��4
����{7·n���(*�DʍLd����CG�r���Î��
�H!%_�����t��������8w���ŕe���W/ou9{G�"��u�*\K�*�xy����s�uto���k�e=.�=�"LT�/�a����9��"+;;wl���'��<�V��X�-��~>��U\7��Ixyz"�0�.]�ԙ���IF5�ܹm3�O�"e��5? ���m4�M�w섥�V`����!���B\N�����ӫ|����7�ǩ��Z��K�*�%�h�kK�b�*��8!�c�Z}�&�a��35r��e�����+�u#M�527EbJ"�NzR3_:uĪM�e�J\����4�aB$(���\�xx"�����kā���wm��#G0����ܦ��lX�-/%��� ;� ������}m�A�s㚕HL��L�;����c�0��K7��\��k�� ��N��G�sԴ����e���=}Fl�s�h���}<U�����w��e���ڗ�����kN��z�EfV�$��\�~��6���s�0y�b8М�Ƕ�q�z�p-๘���^�4!V\H~��زaR�%#'=;֮�U��ƌƟ�d>�"-X�'�d?��G��t�Z[�I�:�/s�#�rS=��_���b_ �6��Oz�_Wj��dt�?v 扞|5���:R遞}3OM��U�π��<
E���g�µ�d��Ñ��4#�r���S���W_C��[Tߴ��֪o��0� :w.��}\����N'N���gn��0a1��?�f�BfF&J*J1s�(������Ԟ���|a2�ӑ�s�<�:	#�[/�[��D���}I�#;'��M������7u��`������ٷs1nT��������Ii&bʴ��}�P:S�M����Ǎ��+'bu�p�g$&^�S�&Qʹ�UUV�䉓�Bcp;'yD��8Y��P��Z�99��Q�G���勗��oj�G��Pq����Ï���qC���*�	˥K(&L��K��1�ʱ��bj2��
sQ����/����#��h����$&<5	�������|���%q0����o������]����/_*���VN6F�y^�>�r����Ϙ�+�ѷ_?q�7.>3�yn�����y�/..>� *i�?#�r�Tp��Ť�S�;<C�h���l�cM�w��"������+ג0��'�(���A�{�O�F�������{R�P^���U�<��t��,r�����SMhW�F<(����v�u�<��V�=�/����xqWp�}z<:cǎA�f��,|J����{tG̩S�4i
�C���^y��TF�G��as�5i^�{�@�P:���)�w!8�.���O�ƃ�h�y�/��*��"�58����"�a#��-TC�L�-0v�8%,������S'0"l$�C�1��o�[�~�0$ğ��BѭG_蠃������g���0+��ب�5e���uп�hߏ�[����.��ܱ܈��8KA�B�Xn�����n�U	v\o-�Xs���/F�_(7j���K������	ڝ��p��5�Ck1�Z�7h�xi~�j���ׯ���X��ߠa��k<�!�R�N-��{�x1���;������q�T����s���4bD����(�7"�uK��r�i}.�4T���ݡ}����~�1T�?Ɛ�˨W�!�Bh�����`�ʀ�����1�4'zQ�^�r�}W��-+�t�_��K���ں�t/B�.��}�K��f��t�oCG�t�G�IwjYt�A����<��t�At�A�>t�Mt�At��_q��C�������� t�At���頃:蠃:�K`(��.N��㇨���9�8�.l���bn��?3��O���_d#� ���u"8���6��^N������ �'[�4����K�"�x>r|=�~+��8j��vp I�����߬.�*㶩���'W���y�1�y�M����x�t��A��8�*nh�ӊ��G���_�U��ס�%��lA����/u|W�����HzU����u���`�&�@"q��3ГH��P56#1y[�/$6�(A�MuK0kh�_MZ���T7���/ί��X�>x���Y �,�B;°T_~�'N�I�;�v���τ�u����~�!��Q[[OOO�{{�m��46�bՏ��w�nAL���#�B9)b|����p%��xh���c�'���E�G��曥8s�*���Ӿ=ޤ~98��Z epT��^~���U��a�*9|YY7�7�������a9�m�
{k+8�8ᅙ����ߢ�7_.�W]Y/�vxy�Kps�lQn���ذal��E},�S��6�_�M�6	r��䄷��k�ƪ�˰+|�XP����3/�D�N���wh���F[ww�����ۢܚV`�Ν"���%^��V˭^�-8 ���Ƙ3��t�ޢ�]O�5�����g�{�]�[�ۺa=6o�,М�~��ԢܪU?`׮�051����{�y��(���<x@d�`�M�>�{�jQn�����F��E��gf>��^�[�o���p��Eeu5��3}���f�JDE�	y�^~�V۷��X��E}�eaڳϠg+�z�F�R��v�"���o�N���J}��@}ij���M�1=��Rn�^1�8�f����R��;�bݺu����{n�Y�ջe}�����E:<�t0�����@�r�����-�Q[^#j�T�oh�����mݺfƴH����'�DG�?��X�Gq����H��D
#�����������/����	���e��Ш���95��x�3�g�WG� �� hf�?��z��A�uvƣa#EZ���!��jki���H'r�h�'�����۶b��]���r���53���'eq"�H�8g��E#�T4>��A�7����ڎ��>Ӭ��� /�s^���3v��ı��ERm%b�G왓X��XZ[bۦ-ص}&N{V�����(+(�[��{{;�oߎ�Ç1a�4�r�ODc����Oalb��{����=x�)��ħNǅ�g�������H�g�lڀ��z_�\$�K	�0g�l89:��v����)S�닎��س��Ï`cg��QQ�i�*���b�r	gcMrx��W����w������fk��z1QG#���`I�w��p�"��p��Z��$���cx��D��j�^"?3f�Ֆ_\,��ěo�&���8L�}'��+��|1�Ob���hG$���HDFjA������D��EP�u�Wa����K�z���D�_���'��(�o�҂�%]�H�ߌE�~R�1�Oc׶--�Q�/��<��3h۶-"���k[���4���1o�;hC��(��ر#�*�8�p�rΝ���/����/_ƪ�oA�r�2�����+��E��sg�7||;he*)���m�>�����>x�]�>pH����"�+��_��s�"�GW������L���gf�۫������c���Z�U���0y������y�F���oQ_���xn�Ӵ��i��|Eč	����D�e�~��s����r	{���ݽzh�..�����t���!33K�~�{���F��Wa�1}�x{�Cl���i<zP�4�u�u�v��=�W�RG��?�M�F����^�L��v���	��X/M:����-��''����*/�����6@��0����ĭ��M������II����R@�n�y�t�B�r�ї���mߧC�HKkQ�")��.�jˀ_�$)Gg3���B���"E�]�vȔ�1*q3�:�-��Rl��o�N�o�6�ȣ�4�U" ��^��C������Ǆf岈�v�O� 񷃓3��o�l��,�����ݫ7/��E9��V@�����O��(-.�����D4��.�ʶ�-�e���=�H�����9"h��"��s�>7��{�}76l�Ԣ>�~��-��4nLO��ͷ�Y�&f��+�UT�]D������ �� �vk�	Z�����%�j[~^v�lY_9]���Sm!��ԉ��i"��S���t�v���s>͝Dj��������ѫ�d��Jd�����3�ł��<_B�ꆝ�CeE%̭4�m�����%�� ��6�7a�[�����D�{����)��bI����qCX���W����KIqq�\�{ˋ�X�����QeeD��P�*�����瓪��UR.Ԧ�*��&sGYI�ȧ:d�Pzƚ���'��@ee�V}�ťHNIƀ�Rߐ�*|��4��r�*�l�ѩSW�񵱵��cQ(.*�������tXA!݄�xQ�I�`#����Fgef���]�����c�:�<��Co�P��T5�5v��Ɩ�)��fz/&�[blQc�=v��wl4�  E�  �����{w`Ib����9�}�������8S�#4$����u��wA��(��?I��:�����r����?q.تj	�a�B�'���&�V[�H���P������Q}��V#�UU].K��߸V���o��5U^[>�rR[k����������i��y�`ӥ+�|�����ލ�^xICn�#i�':]�b�~�*����R_�vD�e�����͛ĩ\�~���~Oww���a��%��5�Z;����p��	X��bۦ-x��W4�:t���sq��!1g�mތa�Ӑ{� �		:u�
�8�g�MxZS��f�ݍ�3'`L�uά��s�hȹ�v�;s�ؐ��؉�FiF�wqv����)�����cxr�x�v��زaS۴����1�����'��q�j\>uB��?���_{U�<{GD������D�����x�E_�ɜM߼��ݾ���fΘ�����O/�\� �m_��~ضqz��Q?;[�u��&��~�j<1J3[�KfjvP�;y�e�|<���������Wwa�l��kW����5�����b����ܥ�<}��Ր�оZ��b��M� mݼ�G�$�&u`-`An>v�|�����KУ{7��r5�5ض~5�?�6m؈��u�(σH~me9����t�X0�'<?Qs^������[7�AG*o���;f��\	|���ho/��	먟�	V%m"L��X��g�1B�=ۺ�Z���ŵ50@�m��m[�`��P'n��pla��G���7~۳=��`� -��g��*'�`۶l���E��^�/�>0'"}��~~t0V.]o:�;9�)�����kU�S�]S��ƞ���Ȣ����`�ܩ�I[-��q��2����P_61�/�V6t��y9AO_%ɰ�S��A����_t6�����^������_��&vrcK%�j�-Y�ڪJ|1u*��h&�bP��T�Y����'�)�B��'b��S�`�ڵDd���{�[oM��v��0��g��9D(,���i��L�������:�ϛK�m��π�?��1y�X�|%
����S�@`/�T8�~0����uk����dvђ2ǧCGL~�M�^�U�x�H���\�1����3{6mP���˯a�(�F�:w�Tޢ�Fs�7r���W���Bn9�GUm�{�E�R��o;an�e�����?m���h<{'W�ot��� a�1���''h�����?�ڥKQ\X�I����LM��ꁗ��˖��_�n��Ͽ��Z�}98���_��=��b�ȑCmQkߡ9��w߈w����א���O?łph�o��S:N�64��*�����>�(&Nz]C����)�͝��X���Ͽ��V��o���~��,УG��R?[|��7���T�ٹc�xc^Дc�Ք/����?�����I��ѐ��s��}�y�g���"�铓^֐�|�o����f�v��}1t�f�/3kQ�'}��txx��Ø��A��7���1�\��������>�"g�7�~/��쉘v���mx���Ł��JY����4��i^���S���s����_�mx�w�j�",�?_�l>/"�=��T��R��/h�t����ZōK}T�W
�o�i���oك �R2�VC��@83�ÿ��	���9lm\`gk+�+��s;{�\�\!���,e%E�)(M(l���ˣM�&�ƴ��ʫ,-��Z؄���*H.��,�5���T���ރq1pqp�jsS���� �-E-b��_[="�v6�ߕ����BҎ�ٙB�U\\[[�\mE���>!&F��365@@@���
Z��T6�X63GiY�|d�RI�5V{�ݻwER��$�[V}3���vV�pn��4���g������Ѵ�/ȃ���2DuY	ͤ&���d"ц(-.��G[Yy�%�W3-��D���ψd9ѷL�RCkt+=�y�(�=��J���"��%X)/�g9��4X^TT���p;'~�d�i�0�$r	1q�26AjYZط�}YMo��t����D��B���WV^Q^6,m�Z�X_>�efd`�c�ZW-�z�&LMq;3N��)4P��(Z�*`ceI��y�O�RJ�"���|()-�[�<@e�W:�#��]�AIq�0��6Kݴɸ�qK\��#���)ߺ�B�[I�⣣QUR#cC��Ѽ�"����;4neps����q��bNs7/� έ],/%9	�.��C�}I��D�������x{7X^d�U����Nn.F��Q��Am]����{	�?��J#�#n�0xQ��� �fL����� K�����jU�[��TS�A���/��&^=�I��[P��k�����&���|���Nb��ع�c���r��AXX�͘)�-X��:�ڕ+��/i��mNǏAХK�q�O�pK-��a�����>w����"�j0~�>S��mڸ��QG�\�;�/4�� !>}�9Ο>��?/İǆ�s���R��3'����c�?{>�"�t�/�7tBB���;���FFB/�"�cG�s���1���1j��9ss����<Oއ3g �@p����i��Y?NG�^����������:H�M��¼9����K���3`l!#G�O���ի�`�B\ǲŋѫwoѶ�o��z�ѩC���~�Lr		Q�9}�8�}o��!�9	�+�O�ȑ����o�����~ưaCq��U|��X�pT�mۼ?̘��IX�|9&�����&�'��z�NP�L�nn��a��9��8�+x��W��)#�Q�WD;R�&'����F!"</Lz	.2_���0q�b�ԯ�\�d1RR���	�<7o�ƺ5k��O�P\TH혇A�ƍxyl��T2bh��m>�y�~{K-Ĩ�T\�~���[p�m�IDƖ�\�o������M6_L�5��c��#�M�&��۶cʔ)D�J1w�ODF��g&>O?��\Bt8V�\�/����ز~2��g��7t0e���0lX�oM~�&�XJ�WR]�3�Oㅗ&���L;����_��~�yUU]�%K���ڛ����)|S⣱c���ƛ������y���Gs���
�̔D̞5��;hab�u�V"7'999�ڻ�����D�N��ؖ-DyD>##"1����[�,>�ڶ���{� |�~Y�@h��G�'�׎�d>�y���L����'����Ԟ�kׄ�<�<�-\� o��&F�~��-C��n��[�>��]��.��bs��/NB�ضu#҉���!ѧc�(����ľ��0j�(���c)�C�Y�gћ/�Ht����A�Aܘ��C_��(g�r�xU��1���Uۨ���V_7ĺy��
M�^]��+ťv⭪*%�_rt3&h������!�>���TVГ���t�4����m�v��rSm�ꋢˍ�sI.�ԉ����<G�~�9������L��ڬ�,�'���5~�3x��Ɉ���i���6F��lt��N��x�LFz:֮]�g����
���w�ٹk��hӜ0AA�Ew���;W7�~�I�ц�|�jL��D��Ni��a��.>'����uk������K��Ν��gvpD"��j�
L�4I����Ʌ��Cpp���B�"�m�6�9BA��ee�V���Fҧ���-�+��� m�%�x�G8���OZR6�YA��i��Jx�������b���x��g�Mގ�OTD4~�u;�v� m�Ғ2�vv��������_w��H�\复����Cpt�g{z�_L��޽���18<�����S|�Vߚ�k�=� m���|���k/�5�f��Q#G)H���B靖���`�߼�<򈂴����Z�6>���ЎHc�.�c���I���ťw�[�4)1A���۷���1**����/o1�ƏKƚ�kh<Fs��jee���	�!װq�V��1��6�ܪ�rq�C��B�އG���2t�Pi�ȟ�U3��� 4N����Uk���_A��e�0jf����	��NĒſ`�a��E�RP\R,���и�����$�u�po�7T�+ R�gl���O�ͭD�n��Wt�ԙ�2�K9�9K�_������è��׮&N9ic��a���?�v�ix-1d�0,^�}z�A@'�qLS{��{���c��������Yَ۴��E�����G���\�Z\�y��ɔǭ��%:����+���e�Ïְ�/k���(j��>�eۿa�_��eF�gm�0���a���(�������]�>���0�������j��^Гu�N�� @=p�*ʡ|5T�t������`�ldfd�7��ŋ͚�WF+}�<�z�8������c>e[[[�ڵ��W�LV^ >�����fD��`���Ν��1J�/oo�����[)L�|[ؿ�?�##In����[��WWW!��m�0Κ��O>�k5;u���u�R���Z� ڼ�B�0����}���?oLM�Q@d%..Vl6gϝ���O)�}uV/����Rdfe"���ᛠ*fA��&,�AYe"��1��A��k��bSc�S��(W.����bD�_��#H�
��b��@�U+0�t����t��&4�BAV���܊�0�;�D���������!n"��R�ny^�`
�"9���돰�P����Y�T�._��K���^hh(� +O�L�B�oz���+X���~��!��E"��`��\�����Ŀ[ڷ��������ٳ3nZ8��׵ �onn�y?~/~�v8P��r(���t}<B�M���l�8^
�,H�5j���l�󼵍5�O���[c#D^�Đ��A�91&\A��~�-�7{&��p�F!nP�CNV[���ө-�,�!22���^EB|4�c�-�ւ�Ξ9-l�hޅ�g���#ǐ�w/��}˖��P{g΀%���(t���qq��$�C�p�~����O��с��"5W�(�&')�ז�Kv5�ᛯ�y���˘@�ݼe����-#�m�|����~?o��ǡ��|�6�V&\�d.ND�9����8ٴ@��(�9&"~d��MЭZb�O3�����X<>�q�<u1��ɉ�����Z�ٵ����x?"֒��HzGe�>ww�&r=绯вEKD]��Vg:X%���>22���.�[�j��l�q�F�x'O��w3R�����:�� AEY_��։��u=�y�9�Ͻ��=
a~��|#�ߕ�c1m�l\����)&M�,N�O��u�)_�6$�\�܋�$����9���N�u��^�,|�Ν�Ƌ
���~rD\l� �/Nz�ֶ��U��߱+���#n$܀��>^y�M�X����s��)ڿ] /Z���$�Z���o�C��\8C�)_e޸�oڂ�������	�G�p�粖d����2ڸ_}u�pT�$�����y��8���/L"���+H��_�`ڌE?��o��6F�S���s��%D�B�V������I�O3V�	r��Æ-[q����7�Y�4u{����18<ʴٳ���ʒ
Lz�5X;8"��i�uv��8"Πv<��x8zz�g�+��sr�ļ��GyY���,��Qċ��j����=pA�Ϣ��?L�Q�0��֢�R#�@�]�f�Ad7�qD�]�X�<ptUj�8<|��TVUᳩ_�>�A�b�ܙ�1s�,!������pv�BLx0���~X�V�ضs7��"�o)'9�� �ώN�rܧ�6n��PQT�'�QyD��i��(����?̘��g΢��� ";�БF-UnxZ[�c񒕸t%%DH��cg���͞<6W�é��E��)_N�� �R{-�)��n��C��*..� "E�1����J;I�ϧ����042B����ꂁ�Q01���m�u�(�S�ޏ�o@ z��*�Pe�a��s�ⅳ�HI���^kD�~��F��T�V�@hHғ����/�]���իlZ�T3ƻo��4��+��p�>��4�Ry.aӶ���e�%xd� x�@`��hV�O�C���di����t�����㗱�m�V�0����+��Lh㪨��%��2�A�fJ�S�qy"y�vv6��N{�_aSل�|E�\=�G"W�J�D>���>�j>��rT+O/K|��?��v���g,��9S�m��QE���2a���cW������%r���j�spt��aRg�v��7iͭl0j�4��}�<^�*����~� ;x��F��L\��jrZ������ �6�����_�~�7��:kșXXk<��������J�����������ghl������Az�O[y���WK&�Ԡ^��{U_C��)}o�����l�U�J�ff���Kչ�MN���nj���\�����:4=������ɡ#n8
���ya��T�I"1�2����^~��zF"����3�kd1�8�w���頃:�Cc�=ڷ��1t���F����%5�}V�[�����J!ǾR�M����F9T���1�**N��)y8E�6�Z�Wb�蠃:���Cc��A!mq{������˚295344�����0��\��\[�8�һG"zΉ*/������q��:��:蠃:<X��L���!C_a���h�݃��+���ʶ�4�+��?�E�����q��焣�:��ڴn���� nl�����ڒ�������`��S=1��ಛ�zЯ�S��426�%��O:�8qsS@���N��bM�ݪ�Ol��To�
RG߲����k�zL7���M��������s�%M�:�"���'�m�Q��o׎�so�v����pFD=Ӏ:������K��j�Q�"���I�r	1�hݺ̭��K���c+���jT.��˙�U^jJlllay���haO���$��յq��X5���Z>Im������=��L�a��ب\VV���x/���3��C.%9&f&ptl<�%g��N�N��dg���.����e破�n��sAN*�����x���A~~�=��+*,@ZZ
�s��K��C幸{�S.�N\=n>�`��<<���,!)))p��mT���[��n��U���p �^���~�����nF
w��fd(����<�[S��tu�,�'H�~����xLxߕ�F���:���9��ޘ��_Qh� ȍŒ�#P�{/���)�B�#b�7[�u�����0p���8�կ��`�A�� �{ￋ��}�G�nP��� ˖/ň�0x�04��^}~�1F�נLme�-^�����'ǣ1L��^��Fkɵ)GuE�.Y�N�1��I���Vb���x|�X�p{��]�v���k8`(���?>z�ꍱ�Dc�ꫯE̫�����:�_�m���_l����@j���iTn�֭"u���jT��o�FwwL��F�l�J���ҒCS�gφ'����4*�k�nя|�I�rk׮��r�׍�mܰY���aΜF�n܀�w���w�(o�:yɚ5��m޴�tp�W;6n\��/a��͍��ع���|�U��[�r��/�~�ʝ<yW/]���s�[K파��\z��ų�p��i|=��~޵}���`�
4�01����E�W����������`�%L�p�Z���~��`Չ4Y��� �[�y����o��P��Дڷ���ZY"*,�Q░�.���vj�(q����ms+��\i�����AR|,Ғ����-;-ͬ�s#�0q���YiHMKFcH��q��""�F�[A~�L�em�Ɛ��F�km���¼�[
��L��n��|�1�ÀF�[iA�
�q���1�gg#�N6M��杔�sʦe�������ܬt*3u��Z�˪��P\xWh#Cei	����,�,�R=��+EA�\;�hyL�㣯��e�F�����"'�˓�񵖈7bahl$�j���UQ^Y)ri�3�n5�ό���"Ȯ������K����cͱBȥ�B�Q9�SV�-ܥy�cآmdb|j�~�4�8d�V�U"9)^̭;ٙ�shXk&4��X��7(�J�eL�z4��KM������ ���U��!m";P�f6��R�ſ������
��S�����;�K�z!��۟=)|����3����zX8U�"��_	����P����^��Fé�BC�hm�1�����Kx�} �cb�H._�#"�]�O?�V�[#::9D�����aeaI�E4��D�utp��)iDn���	c#8�	�Mf��T?''��K2h<7�:���VFF�r�Qhne���B�$�jı�#,�**h��KMN����V�+A������pP]m����4���N��%N���"ppUU� �^Z�w��w%�E( �����u�U����6k�	QQ�j�=~��w��f�	A-��7��Ef3s�;�}�F��BDsֈp�wמ�]
bhޱ9�MmgN�D?-�Qa�d7��E�.��Bc��8��9zG�4pJ���5�h�:4u������o$&����4W�����&�~i�����j��#!��b`�̂�Y8�5@����f�ZZ��^���j���ȥw����m�d�� qˣy�G�>WWW;t�{M���Z�y��{�:m[��_I��K��ɍ,H�&F��y'�:�w�/�_�*������Ik�^��rB�i��h��F��}EB��"(��t��;kW�A:
��[R\��("
�k�	�ܱ���͝�����[b�����i#f��^$��z!�<=�wlGVfV��-6>F�SSSӐx#�ݴ��{��'� �b���"n�qx���ʦ��ֻ����F !>�6����[�V(����chr�D�yd �*+���� q�THCD�;Y��l����LF玁�x�'�6H�.]���O���23�$n�1Q�գ���#�TCč	���O�ƍ4��$n7h�z�z���|�R�č#��5׮^���L4��D�m�$P��6Dܸφ*�Kƭ��c����#z�鋨���"P�;qӣ�F6H�n�'���}��A����[Td$�w�"|~�C�$ni7o���+�t�Ns,R#P��	�x�vv�l�4�����B�]k���I�Ѯ:t}�⣢�%�\���Pw���8O���+�<��vM��K��_�q���o�4d� rl��Nv�Sߍ��D�1�i��`I�!��߇�����{5+-�y�9�EeU%��B����,��[Ϟ"�RxH�Hף>���ͷ�_�&r������]�u� "ϝ�>�6Ð�P��l2Μ8A$.���f;ؤ�Įc�N�HO��"���q���+W�fsΟ'��SC�Mb��W�~����B�榴� �O����kL�������\��#������F�8s�֌���x��_��6�$�_�CGk��kI�:��/�~#��sg�_���k+��]�s���}K�߼��O��wD_|��Dz3p��E4��ǎ�	aM�}���8T����}��B��w�������8���OO�}K�X�CF������S'�����۶������6t�Z�¢1|�6�Z;~/����iŲe�7��Ǥ�_����lX����ۏ��z-��o�ְ�٥KAx�I�r��_��������KA��(x���1}���s�屦���GD.�g�hМ���੧�F[//,Z4�СI�����]����Ӿ�O��p�	u������c���_�n�n�������v��卟f�BNf*�4/o?t�G�D[/l۽]���4��o?t��0�ΞG!��V����{P]]+4n�����޽�:�+0�u��q{�/TW�;��&1�#Z�?r�T�]NPEEY9�Qah��R�Ŵ��p��-9�P�� 2֙50�f��o >��}<Ɏ�j�\Dx(l�7���+�s�����8w�4z	��!�����h�ߍ�hX��Ǝ�s��K�Od�F�,?ӳ��x��}/�:Y�T��>���;�����P���������Ʀ�����ƍk���<���_����0ߺ��c�� "l��gu�-�\@{�޶�D���̴1�B�[yY���i�_hH0��k��Y�a�ʕZ���~�Y5��K�5���l"͹4�-$r�D૪������֘���&�*�ˑ���mag�&�&���BI~,l���*n9r�"sK")6�R�[*�GK{{�	tl儸�XqH���n��ɉH�����Q�#;%	n�ۑ��q��6�j��.���,3%NnRmibL� �~�̛�"+5��Szk4;5	��������0u
��E�PUd�'#>6��LTV�����Qa�n'�Z��&�dʭZ9��N�����T;�p���׮��SQSS� �gZR\<�������ik-r�&�LDrb�ȷ�����]:u�(n>?���q��TӪfg�"62��{�4��#�F"����Ң<�J�[���wtE�֭���s����6!2C���;q�J��Yč}%����Bk������kA��G���$�A1��o`ng33D����Pi��?�r:T��=��y}�+"T�t���*��_ն�/�i
ȴn�en��3�U�UʋLS >.�N�����������AZ�M���K�\�k�]�-�l�G''��]��������	���#33�Am$�I-��DL¯]�9ٷok��Ο;��_=sy�yHI������M��F��$�'��]�4���ݻѡ}Qy��3�s��E"��T��7+*�|�2m�y$w[�8�H�TF]��W[O\8u������u"�]%�(��y�RSSq��)៓�{G�\���A�Ù����/�Fa!���[U�X�Ąx���	9�8����ƍ8tU���`��O��,�����k��d_�*"�OAYI9
��&��A�N�<.��ؿ��fp#�t�6R�<�l�kN$������2nј�i��4^-Z�	"������왓5n�D.��acc��G	SnuM%���Չ[tT�Д��fΉ杝�q��E�U#n��E��s'���srr�-��jč}�J�Jz�
����!��:q�N�1a<y����ƆF�<�>��bbp� W/]�����Hu�E䩕Sk����x[X�Qߟ��j�-��sbR��5�"Rn����5޷�g�����S�`ll
#}\�C�:q���R�ݻ��:5KJ�C�� ��č������K�j#c��N�R�S���Bk@
�\���{y�J�� �׮�yB���t�P'n�����$�ĊKA���9l
0ᮩ��s�hB��o��䤗��W��x�����*!�kD�^BaB��֨���z�������A#W�e�v��z(�]WU#2ẖ̌�8n�Ȕ@��c����N&���4��g�z'U�R�U�?�70�5]��Y+&�����W���7����O=���>2��ccmS����E�t{��������GF^��,"wKQQY�s�`jl��>~8{�<�NT�ڊ
\��.ݺ�&sR�����s��F������X8�l�c���X;!��h�O�9����q��챰���?�~ʍ3;�}�B�H坺p���h��Is���∨����M��ȯ��� ��*�
��N}`F����������+/J�[]e)��Ex{y�ı�prl�#:>FB�j+�'�����������gΟ�7֬ݼq��&8�� ��۠���(��ׇ��,CPP\\]��\ߵ��^�����[�\�_�xX�X���b����&��A�.�=K[k�І̄�ۇ	�Iy|�4/��~����dM���j
������S��fV�pn�,|$�V
r��AII	�"F��q�5W�زe<=<p��"F�0��FDL<V+{� �1Dܚ�[�AC�/-�����fZ�����,���Ҳ�b�c0\�J�斸rF��o<Dr�۾g������������n 	D2$�nk+�̅���+p���������_��A�����7SD�Hcܺ��WM%Zd��њ�}�"��8s�$�M��C��޾nee��� �T��EE�%P�{Q?_�zUd�qw�sw���Bu�O��`�cek3�qq4���Zy9NP]<�<p���ͽ�0=OT�u�|#���i��p#�o��!��<�U������+��_D�F����B1|�T�Ϡ��F&f���M�&s��a�C�4�_�aj!V�Z�{�5^�\�N�Ǯ���z�CղO�M[��+��_Ag�'n:4���B����s��F-Cߠiho����>�$�ZѾR��{��*��a�D�-���}�%̛7���J�����J���ޭML�8������!�6���w`�Q4(��:.6��a��0���U8rp?BB�1�6:���.�N��^>x��w�к53i�'"�{�.��b�fV:��/_�2Z�͈�]<{�v�l\���=��]۠��牰:tC��Pl�YYY��`���046f� z���K�
�?y;����sp���~���S�q��	��S�daX{�ݿ����'�Ǝ��%�������j���{p�����w�ލ�w�R�P�F��l����1���~��{��"
�fnvFO���3~�*�[}D�7o�(ȳ���2�?��3�l�*"0�У�Е0k�L	�`G֨���l�&"�G����X�d
r�`�Bf�䲙p����D�e���pL�r�乬�9G��ܹDB��)1T�ʕˑ��{g������/�.$�<��~�}�^y�u�Y���lZ�H��~�4����ϓ�U�I9=햐������租|$�����4��\?C:8�m�/�|*1��i�����>�u�f5nRy_~����:����&��'�~���=�������+.���M��o�nGM���x�7���*�}�'�ZB��v����UB{���K��,����g��ܵD�����{��Uj��>|}�	�u{L���o�O>�e�a��6��~<��3�޽� ~�1�0���88���1����R_q�����Q��߳������� ~$51^�d�i땇�˗������4/Mi>ec�g#���|d�(�t�4������ ����J"�����3'_������!���wI�r�s���s�z?+"
~���s7k����֩kg8�)�p��ɹå��**,����*�/��t�>{�r��*�á�vX���-m��Y�iU.�D9X-43K��%�`l�w��R�)�����z�0���}�a�/K���;�z��!C������C��6�LM�D���(x{��ݧ�v#=���!X�j-�K��+,*F�=%�q����۷�,�-ϛ7Sac�B�����5`�.YN�M��J�ҫO��'�.�np��$r��h�"x���)��k��X�l���}�f�n��;8�@�U�{G�W�^Y�֭��;��]��]�016���W��������h���X����.y.��m�l%~[�TW�f�Ȼ�� nii����Ak��[�4�:t�k[1��:*�K��V2�&�����[��VZ�b^�	ث�7���E�qy[�ۣ��}��9??�ml��+��Ж�����U>�n�ξ%\=<�ף���X�������&ݸSSt��ӳ}�����_����<';V4W�z��	��0	sqqCe�Ҕ��q#w&h$D�/�v�ޝ�얂���Jk�&ի׆98���m[1��ro�ѡ:v�К�xx�����Mĭ�_r�P\T��N��:&u<�Rh���-�HZz�����C388:�O����΁\�������e�BdQ����N�e���Tżg�lhl���;+�N"CKAA>t�AG��c�#f�򓟞����!MA�}�%a�T����J�����"Z�`����\)��G�E��V������[�m��������D�ţ-�y���r�>�`bj��\w|��4�VI���=�!xA�N��N��c?*U09Z�x1�6e(���Ǡ��L"Ǳپ�66J2�YJJ�$r���y��֊���聮ݤ>=&�V�>c�$��������Y}��q��G�ܰQ����TLMVv�3o����yt0zh����̟f���N�gr�ةTMaf�/�gσ��R���=�@Io�:嫩�F�������E=����ϦP?�R|���C��$�v��7�%b��;����F:�EK�iT�_?"�?/\(�����{�K_"l}��F�ܯ�.����׬��{�}L󫥲�ܖT?��9����V9_�v��H�$���ާy�4�������?׸���_��N�Ϯt���o�����7��x�v����)��`|�ѧ"�<���k5��>�~�C��U)�q��Ŵ3��I/0Mx�Y�P��>���ג�<�q�˯H��ޘ��
�&ǫ�'��Fi�w��i?j�q|�I05k��ES���<��<t�*��¬�a}zI�Z�o�q�ᯅ�z�'G�"��̤��i����n�=Ι�Z�K�FNnj�E�Gbחl���z���������"�8�P�^��JQ"#�Z�$��6ڄ,�V�1�P�~��u,�m�q�?N[�����fnW[�L����W%m�
k�C�xy����������1��x�]9��K+[;9���4f�V�>�H��w�jK���Ps��i}�����xܬ[h��f=�� ��ch��#���\'���Hl�eh���E#"�즙Vۼ���W[{�,��5F� �{n���p���#n�!܏�M_��q��2����.M�:��`B�^Z�'}a�mV�����bk�kd�I�:7� ��Y�!�ß/:��:(�gͥ:�v�=�Ǆ�^�#n�a���j��{��o.UU����F�Aח:��_�o�����i!��=��M�q�	�Q�`�i�Ui}5y�R9����jj�a�g�p�����Օ⿪���yO��=�M��&����l_������/9������CC�V�z��O��b��ր���8ꠃ:�~�s��:�E#�{��KCT[�5�W���}Aa����+��2�|��S�B�f���N��>��Mt�A���3�+�:���C�P{̇z�l:4t�:�[t��\�7�4D�^��P[��j���ǷR�U��B�ť�����E01oFT�Hye���&
Ez͗���P��r׭��8=���,����%T��� F�ƜH �&��֏ۢ�9����f"�����"��Z]I�P�*+�9����q�k�5$��ꚆS�PT�W�� �f&��`��aX��F�1&Ʀ����+�(���q}q�Ý0*KK�t�cѐy�%y"��$E��gW�wKXZ����\ey��#�ج��ļ����Ĵ��q��`����F独�4�kjeE5:�ղ���]C�9P[[C"�$�mh`�vT�W�\����O6z�7jx|�X\[Y.�}-��Ʒ5*����*�PY]���ע�\�Q[�ۉ�P6<��*h������p;:���M1#�5��.�ۿ�_���}�D�����&l���bnV�����9_��Y`�c#��
ꑓ�����J�373������4�gRؼe��<�
���
�zTUE�l,�7_,�4~ֶv:l���ڰvJKJ����=����6 o s~�)��33���Q��b�q��X�yw�`bb''4�>����,,]�wH����ha��Cgi ���|�
��������}����rE$���T7��٣g�^��C�ܞ���Y�PN$��kaa���Gk���ع�Wܸ�##}XY۠o���Q^)�ϙ#���yC�?���\�֍������2ص�G�Ν�g���Y3Q\"��ߌ�7�Ʒswi �
"�i��Ry�/ͭ���#�cL�������C+���ԥs}nV%���_�ׯ_�9�F&Fx��i@�4Gӿ��UU�W�����]{I>�����+D����S��Tk��5�V�v�m�������;���aR1"O�֯G'g�������{=��:6�_���"���_:w��CԒ��sׯ]���4��c�o�A��h֏��}�f�����7?_xxxb�Б��D��-��s<������Aض~-"�#ajl*ƥ+�qo-�`邹��}[�������|�&UK�� �Z�ӻ����[�`���Z�@�5���к�� ��&U�� �s&�����.nn9�i4%t�D�Y(��E���\�u��բ#n:�n��@�2�,���H�Ҧ� VV��o���%�6J�82~��=EBnN�Ή�7�F?��"��V�V�DpA	}C��Da֌�X��WIy4s?����Hr�q�:|��4I�w{'g�`�h��ё��z�X�q�D��AB���S:ѳ�"��5,^���0]����|�Q��FlJ�3!.?᛿`���p��#F���Jl8q11�?w6V�Y+�@p�={�FEE��H�N�l�M���T��rT�>}��n�]�ٷ@hH0>��#?wI�/�eA�4�6D}ڰ������s1{�|�[+��s;8珞��������q��IV	�k�޽QE����P��Z�`>�M�%	f����q�C���H�y3g�@����,
�<d0J��!"���`VI{9(r��=Q\\$�-ݸ�/>��v���:��|�EGG�]W78�(��r��]�����\�S>��7n��J�ڎ$�^Z\(�.%%�Y��n����&�I�q;+�(R�����GRy�)��,R1�߹#TjJV�\)�/8���؅����"Ht*�ߏ�+}�4�>D�ď���t6��͛www�@�z�޽�����sJ�)�}�_�,�F��ݺ����А��c�����8������'�7N��j�*�{zh�q�9o__��ȼ��y.,�[I�.�8h� �t�+�+���+��ڪn�щ�iKG������;�K_��HϞ}p�FF��߹8~�8�Z�c7U�j/o1W*��[�d	<==�Ou��q{��]�f�V�o��g(Yh�鴻f�
M9j_�>J����V�X���;�j�����ݔ<��ׯ[�5 �k��}112r�Y����F��M�ؾCJ�P�
���桼�D#�@@��;99��jj4g�j�8�8�������jd�P�k���=-34�[Oe�h#;v�$���*�0�ϸ{�Nde݂�
qS�_��g�.�?e�J9��Q�������ӧ�P�ՈB�Z=�f�Cn܏�DXԉ[G������ϝAޝ��^�nD~ݺ%D�ԉ��<� "����E�_�}`�NXBd;��:q�����<DE\'"���������D���h���PiGiA.�b��$I�����/��f��_D�t���2���|"��9$�x���`�|�_!���b�Ƙ��\�U'd���I؁�{���!'�>W���Ew5s�z�u9�=�B�/���z�?����W.!%9Q���J~��q��̀T�����A/ =햎���G5�:�ßk����ؼ�y�*\�v�D�jj�h��U�V96S�Z�A�.���@�I�����Au�ʽl�[�`���``T'N�l�4�F����/��1���Ʌ����m���*9k+1�,�x#�VI�}��-,�y	������ԩ�T�*��5JK�ann*�~��3�[$&�@EY9��-ЊN������u�p��~�Us+�������I��K��⅋(,*� �e�����c��Ţ~&$SC���Us���v*�رi=���e�[7o33s��s�ml$�mX�
AAE��/W��hf%)o���8r��U222���**��� i����q��E�K�o���V%��ܝ[��܅f͚	-��155����y�
�:q\<����?����=[�c�}�y�ҡ%r�䡼�R"�i�*�<qB<O^G�cC��ٻ�W�������~��������氙e34onS5���b�͢��͕��a|3�ܹy:(r�ѳ��L�:`��_��{����v�T���J����mt �Mhh��`����4w�};q��A�3z�ld�>3+��JM�O��_~s�����+���UKgw�����c?=��5�q�ӷ�T��QlذF�>��˃������I���;K�*;;K��%�GNn�?"5!_�xK�"L��ƔW�������&�s'� �K.v���'��e����SQ��P[�L��X��ö���=)+C���Г/�i�A/  �*IDAT��~�o���rl����vGS��W>x5�,��FߠN�j*b���Ko"ڦox>
�"�O��j@m�pRV�xJ��p���V�ZXM�/�~��I]S���s9����0j�T\ΝAZF^y�uXYY	By�d���������«o�*6K~��� d���@�|��ჴi���oO�~��@!��h#]))/��bRb�y�=TTU��+.6�#�QS�|���څ��[T�ɴʒ���Db���h��'��t1��S>�t��o���#.>�Z��C{w :*
o�������B�$�ڵz*/��9����{TѦϛ���l�ؾ�Ȋ���ϝ���`�6�Ad��͛6R(��z�*�.^��$����a&y��F%���ӧp��e����0!2dbd��	طg7�C��E_���{��_
��bZj*��e_�Xէ���˗���W_�%�����x�o����!��E�!R9�ɧ���-L�9�s��O?�Q&�O��Þ=�0��7�˟�Dҙ@���1�C��w�Es�L`�?l�_��J����ظq�ho�L����P�了*�#)6�Ť������ɹ�����5e���Gc� 5@ʿ%��Ïi�5'"m���xj�Iaޗ#9.
�O��KT�_��R�|�r��aF���8,[�o��6Z9�F%�/�v6��<P��a�#��`��'�֫� 0y�6�(��ө~���ǟ
��ĸ��.�.Y��A��w�c�gW�p�|��ג�䬍�?o>�|
���4-����_�l�*��wlێ�	.��4�};�֬�ȱ�t����k����Q�sVf&6�_#B���`���o�N����v��#)��� �n�s�=O��V()����PY��ٙ)XO$p�SO���A��b�ƍ�0�Z���w`��G�渼�\x}Q�?�:��׉}�N�3�>�z]IF��k����˯�R�"^�=K��n���<�W[�ף������g���Ina?O���0i��:=�r���������dS�\&5��.Y0��z��l����o(��҇��P�.[&�˹}�6BktWq���D8�C#�w��ԫO/��:kz*+���cb����I����0�رN��]$���X�v������d�����,-q����eW��;�h׾��TeI�k	��U��k@��KBt8Z�t������/���]{)�ggg'�o��bbhC�@���Ϝv����}�%��Ytѓ�מ6�-�7�\�P��6|(:��~�-�����B�S.]�|��W5!;89����F�ܛI�����P���hj�=
�(����������h��gϞZ&9��o�ͫޏ<��i⻬�D��o!��������Cij�NK�"�����[������V|gm�N�KZĕ;��<��O��a36W�F&7<;v��������#H��wrsy�7Xyq����$�wXΞ�6d�H��em%��:Uz9Rnޤ~����d�ĦrO7ب��Φ�5on��C�I�8����̗[��~4WQ���ԚH�!�r��<������ �/l�3{����0?�h~��y%�wO/\����|����j�ƎS��h�cG���K�R��vx��ae��C~7���:�It��ъ~�,-ĩ��%D���_H4h��~�mg���:���@��7$�_`2y�ap������KBKM���F�*Z9q�W����{4[��5��CXC)�{vE%/�������B�	�bG'�DEb��ݒM����)Hڕg��%�%�y�&n�r9:v���ack�Vtr���ľ�{e!<T���F8F_�p���<{�셋�-�e
�¾��¾�=<<�
���}{�i���T���׮\���ŋͧ�e˖���F,��x�h׾�^�����`.n­_����*n����s��A�+�{Cdfdb��5�\U]�$
��DM���#���+,����ſys�i�m۶������'�{+���"r�E��jUN��/W�q��X�\���~숭J�||�s�tq{���I7n����D`oJ��M�ee�8w���"�;vle�p$��m덣Ǐ	96�1�ٵc��74R1E�)516r�4�YY�ؾm���us%�`���k�8s�x���6�Z�B�i\�������_#4���-�������RU�V�֭��~G�;"|���C�f����ԑ�c}6�ٓ��~���%�1���|�`�anN�;"Ʋ�J9�D�Y�y���L.������,!�v-Z������S&"��؂�W%P��;&�����i���b�ݽ1����
�w�6�N��3k�X���^��I����Q�سk;���8l�:��Da�0��N[7�ٷ�橣���Ǆ+��
Q���������'���!��ı��O��.ݕ����b>����mH��w����Ǡǔ�T���q+#�Ϟ~�wm��#"�I�֊Ɗ/!=t@������ɓ���7K���N��>��>���}{��9����U�G��Q+n��ܤ�͛�B�<PϚ���F�����2'<i�X{P������,$'Lz��� K-��5T%q���|���4
V�-�EEE§���'#,8X"�~&��C�r�
�A`�X:m���9�S����Oh�֬^��zS��ؗM=z���PB�$o��<�,�oaQ��8TATd:�ԔTqsn��tYk�^�[�ވ��!Ҵ2?�q� %���6���z�Ja��M뉱O��#n�)�t��Q#���%rf �|/��2B��`�ByA�5"�5ڷw�ؠX[��+�!8��0�ʗ�n��R��j�2�PYE�%xf�ӈ���Ck�?!_r����gID����w��ce��v�ĉ�b�ƍ������'��Sk'�K��?_�xtP46�ۀ�"4����/</̻�FJ_.vT���޹K�����`̘ǉ@8�Lş0����Q�Dyr?�	'",<L���ċ/�H�x� PLP�<�6nQ/??����V ����4d��id���Ч__ꇣ��ق��=����Z����7�xk�P�f�"9#��lF�� ����P1+W,$���C���#,,��urk�O>�+�-�yd+n��yb,���WP8'�N��o�~p���am��^{��>\ՕUU�Ϯ�ʫ	�x��k�b��%0�C ������D���h�-m�ͷ������$�ǠA����FR��'����w v�U�?����3)��{	���D�tŵ�����}[t�k[{Y]AE�
��J/!�@H!��2�>s�{�w~�罓!$��k��y��>���S��_� s%t/D8CGS=H#H}�{�{�Rv�u��ˌ<�/;�5|Ğ ��3�����}�_-�E�/���9W�r�%3�я���š*�-���IS���){h��۟�����_�1=���<�Lkjh��3�TT5�[�~p��s�=�f��E���ެh�C+q��������a��r���^%���0�&�0p{�&�Nʞ?��}h�e�����-Ed�=��^ʻ&*5��5�@ܮ|��������u���W}��zn�s���������w���l�P��+ߥ����Q��\QP������Է켽>����]?���3�y�so��W�`�Z������\�p���w��ߥ��e�'?�e�]����w����{�����w]eo��X�λ�-�\��Af��z>����}.�����ݻ\���ہK��8�|�����A��{��ŧځ
<b/�Ks�`���
���&���c�_b�9~��cM>]>����\���=f�}�E|n�����%&w��.�+�}�C/Ed,=�=ԸXVN2�r� {+B�d��Z"���e���e)o�C���w��"_�����z��)h���
�����4�8��:\���[y-ε�%�	?W��1.�^^�2�Uz��܇��k\p@L���k����H �}��>���o�u#ʬ�m�UF��<��^��l>o�	��VWTJ%|p�$�n�\�GH�*d�����T?���J$d:Yam�q�p��tɏ����R�J�8��$SQ�ϴ[�?S}6��_U���yR5e{z�[TUS+��|���DG������(ʫ�����̕�����K�Q��j	�,b~ �tv�Ǎ�Q�DIQ�~o������jW]�u���g0?`�D[���kUU5ޅ>Q)�%3f�jO$N�dl������I�$l�����{@�Q�O1�g�=!5X��4R����\����m�U���������4_���pcu�hy߱@�@�������i�y��D���)�cV��b��wI�����i��N2v�B����5B=���I�	)���_�MuC��G}�X�w��y���X#��������:�P�������b�,�z)_��P��_���w�{�͸��!8�zxW��	�#uW��O�2�{�~(��πt�Rm���ջ�:�v�����:�E�A�J�o�CM����+;���ޓ�������d:�s��:|?�
�T,嵶��u�|$}�zzE8�� {�5SU_���9KWh��9IFiԪE�G;z���_��$���?���!��+◺��pFTp^ds{ΈL����ϲo���L�GJ�����T�k_�03���%��CF(����M�K��w�9��&�k�>( '�I���}��O,�F-E��'��2y�-sΘ�{=���_<�{=�2`۟�[22���������&l��� %�=W�7P:h���@�1�}2��_�㾴s��2wV�J�f��� �o!�1+�l��TU��	��	�x��~`
��A]� �J���F�4Dp��R� C�-Y#�~����Mֽ{���z��G�p������]ÿ�4Y>@>XyQ���A])��b�_B� ��t����A_��>�9�.؈��l��U;�,�N U<V) �Єp�!�O��K ��u����1��?��?9E��$x?	?&���^~ \�
�2�JW&$� ?����Y��ݙ���QU["=�N����LF�� ��&s��) ��`�z �:X,��4�eD>Ϣ�2h��"?6�O܂�$�&�0���;�ʥ�0d<�*��ژt����i��T�]��鸂�mq�|V�\,_��\ �4��&+���6��_.�r�(BdYe���_@�uɮ� @dN*��=�U���~O@Iwg��zoc�u�T
���SQ]�v* ]���W�0t���� ,�xW?t���ɒS4��en�R�r�3n����>f�Iƣ|)a=��k,˨��fا �eY�\�*R�k|������Qm�٩q�r��c��i���N�?�,Ux ^ �8�φ�N�<˸�g����YĞ� �r���	q�UD� @.��}�W�:ot��C~��յ�w�b��gOg��m m �t:\�R�6߁~��hS�b�,�眙X�=����C >�XS~؊�J�#����#���Rd� S)�LE�R*�q�&qo��?�����v����L)�(N���@Sʡ��H�$��Ҡ����� ��X�o�iHb��W��#��7�|^ʿ;@ǁ������1���@�=��"���GQ��y$���mTH��X{����Q9/g zq6����ۿ�;�2o�_Y!MB�pH��/mAum��H��%	�$����3��J��,�ʕ����B��� �+/)�X�F�z�n)9v>J�N�B��!�F�Ir��D{��"SiE?��r�A	�;�����d���m %�O
p��.Ԧ�t�u�I�D��ےB<�m�v�T� r1��t����� ��Ms�����~���>*ep�X��a̯�GZ�ʊt�����'$a�f���JH����ch�/�|/�;Kj���eI�ra�Ka�n�I2 �tU��Xr��@�sPnQ �1οEL3ά�)��`��G�H)i�"�%�J,hV�hS�}�	�h�i�Ɍ�RXO�%���K%y����Mh=���EeM8 ���,@�<�y��i\�1i1Y+���-h_Ģ�Ƙƣ�a�����ش���U)(��*[�\�A�@m�E��]Rj��t�h���}���(|�2rr��{zH90*j\+-���e(�����ξ&��]����|��c�}e|=,����ږ��d�g*�t���Oc_��ii=��6p���N��S�����%b{�D� ����_ʁ���~�/�����P��(`�Y.�e9�w)���^4��=��G_�RE��^����$�F�pWD�d���:�F�S�5n�a��L�V +-Ϭ�];w6�|N�:$lF�/�`�T	���� '2��+rIʄ���$W=��L\���##B��/�x�F$!�l�h��ڀ��qE��5[���7�[-/hȍ�vc¤�.�3��x��ֶ;��I��:��G�tp�M<��׭^#0�&���̴i3dn�	 ��zo{[���sD�=VQ� ��M��m��M��@+�$҃�O�-�6n��;�韊vp4dX���z�Zeb,wl��?ۼi�eG�iM�c��`�|@'�k�N�q����<̆�21��p!��ÏL�Nps2d�h	q �L�;[�	� d4F👪�EAb2k%��ϊ_�����1!R��Y�����U�2��qc'�nM� ���c�۹z��Sd2��>�q��AxE�v��lذn ��ƦF�k& �ƥ���yc�(\���2@�j|�B�u�6q�і�g��;��9z\�d�>ȻP��鶭>��DŃ�S]C����Ȝݯ5Ӻc�Ȩ)�5�MS�h� ����m��Mz�9��-�36���;E��!�p�ܡ�b�m�m�c���)fH�F��y�܀�Y��q��/c�����k�5�z��>�M2A�+|o���[N�
����mڸQ�5�����&YӰa�H$#Mc��v���5�7��`�F��r�@r��M�o |�z� ��z�z��sk�m۲U��4�T�G���}/��D�Pؾ^p��
!·}%R?X����"~
�s#�a����;d��(�\���r��=������ف6q� ���7�l����4r��m��9~��7���nw�y��z*m�6q�;�M��ٳ��&����R�
n�흝6����o<�fΚ|��V������aY��0o `����m�Q�V,m7�p��y����0irAs���QG�7��>���_�on���þ�߉�
n�+�x��[�H浴��a�'#����j�����y��>bn�\N����f�뎻5J~��B��sϷc�Y4 >���s�?{�Lh��0��;���-oU"q����_�:�w�n��$��c�/=CZE���+���ÆhD�����s�@�)�>&��{�Hc>Rޗ��;���k<&��'�_��556��
�ȫ����utЦ9���n���Ꮼ����լy;��S�4��t\w�w�/їd<i���2[t�bi4��]w�!~7�����N?�t;��eZ� ��yX	�Ǐo7m���Ǚg.������:�{=ƅ�B�UĒ���ig����W>��}��_�Ꚍ����l0���zz�痵'W��/}��G���C0x��w�ҥ'ht��~|�+_�5<Q�;�m���3�<Ӗ�s��es���?.>@�i���O������'�qDrZ�n�}�ӟ�?I�6(g�"M��O�]k�����	(�.��";ᤥf�����/�C�=׾�MD��˲��ѥ����������/�#g-;�ο(D|��U�o��1:_J����u��v�.��۶y���׾�����s��~/=�d;�쳥ed-����}ކi�Y@��l��c������;S&O����w���4�3�"�[�A��M��o�Ⱦ�v�ء]>_��.��'-�I��J��/������ �jD1�Z����ʋ*:�|�TF���v�y�������/h�r�������w�
����\\=,�no�N<I|N|'�7�;���7�i���� ï����o�����"�:L������h���>f�*޺e�͚9ӎ_�X7�v��чW�����'�Mf�B1/�Ƥ�pPy���Ɵُ~x�֬�*%M��#�� �����f?��z�8y�5�lѦ	�����	$��ͷ�ڮ��;")m$�#~U~��3{�]��~;Y�����߻�>2~�55�����cG��� ;/�0|��_�Y��LUq��C���K߬�R�vAXz�������΁��'BA�W����z�]}�k_��S�K{�I?B��|�C��-�]���}��߱���kj%���3z���}W�WѾ/~��ܫ�T������Gdz��w��־��o۰�ý��2u�F�n]r�4rh�H|�����6��͇̭.�E��� �;�/��5��z1=����o��Bi����{�}���l��"f-�?�`�z��E`�����U}�'N��,��ٰ�ü}{}��^ဖ�ӧ����k ����ڡ�^H�!��4mz07��	�]��F��6_��8����c�i�̕ɥ/��RO���w�a���7l�6i�4����@�Moz�ڇ�]��:��׿��M����
1�^vٛ�q���������׽3lҌ�R���|�6_ϤrB����l~I<ih�	$B��q!�c�Ѓ��}]���N�6S��/���.<p�q�}?���6����ǩ�p�%}�\rɥ�Vd>��㙳f��y��y����?	DQ֮Y��}�ƌg�,���<o<�<_�u&A������v���Җr9b��=���\��6oTʫ�S����X�A>Npڝ*�n|�HA�>��N:�ސxa��_�_��'^���Ú7�U�.��G����۫X^�����]�����{������r��SU|�7�xR��L�B�>�
3��~p���7��H4h�?�lvA?q�l9_c^����k��|㐡��T;��=w�@��!����o�֭�l��)VQ�`-[lD�H�b
75���>��a�vn@���p�9�� F���c�ڛ�y���kdj�?	d��0�����?k---.\�42�� '�2m�%+�_�eg�fW_�A(�d
%�%��q�v�v�E{���]`����%eVi�v>s���H�=F ��γv?Ly�b��z���ʦ���L��:��ꑇvp�њG�T�.P�u�8c��#F��/,������q�>�u 3��V��.[�x��{ｶ�����zŘ��e�ԙ�۹[���������Li�ƌ���Б����VmX����%����9����+�XL�1}��̱_�x�mٲI@���B���:�ڌ�p���ʢ�e�fo�t�u����X͛������A.҉�Ȕr����J$�俇O��nt���m��w��n̌�1Ĕɚ&�C.��Ϯpc�\�S_������:ظ�/-۶lѺd\0͢����n�.e\�X�����6c������������/۶m�|�iґ�w��W�8DcPuj���W�zR�I@K��o���������mּ��ĔΞ�怏K�r�6]�~��+���r!��Hߗ��4����?"
�� �'����ĉ�m���	 ~�BV&ML�\+*�)&p
Q��M-�<Hk��55��|9r�@�ѣ5~k�Ej�R^�\�fΞ�x}f��푇�����M P��� І��qP�K|�=w��|��w���ׁ;��y;(�a�).1	]@�.�ȴQ��0���kXʎ��Ǣ|i����}�WX�#ɿ�p���pT)��=����d���z��j@��q�ߋ��AA�48[;�;f���R/��<LG�� ��^USeu�:i�B)����i�.� ���B�(��H�+�ɍz[[��B
zp����k̘��苤|��U
(�s����뤉�����hZ��M���%�;|����]��H׾>���:�w������MR��mD��45E~/rGWd_�ǨR�"E�3���s����yI��E���	�����mw���G 2)��:l �`�_��];eJ�S')�0R�YEДTW��G�X.M�4��0�R��*������G�����L�[�m8�;hu��� 3��hk0F�s�]�}�E 	�D��r�'h%ۣhJ ���E#����7��&Q�&��� ���uk����5�k
O�@�S�'p�"j��_(j�P���	4�|l�K��ڥD�hm᳆I-��a����.+�iȿ�(�k��/�!��5���n۶n��1�1���u�*� ��r^V.:�T��gGWWXJ'W�/Q��C`�� 0S�z4km�%��A6I� ����@���g��y��F��ZD&�j��ş��:}/u�L-�E�Ł0cX���m޼Ŏ:���������J_���s/ǯ�ou�b߫�q�/�q��S8'c���/S�n�R����uc����RT��o����V�M��L�LC7�����K�Z�_7`�4��}v�oo�c>����SN9�fΚ��E@͓O<n7���L �Gy�.��2?�\(������N��W7
�p��s�=6m�4i�B�~Z��g7=c?�����M��7�ʮ|���dFH+іޏ�O�Q}�^���>��Qc	�Pth��=����G�y�ͷ��N;��]ѭ> ���ȍ�������&N��&G����CN���~�s��L�\t�!1;~��#�ҭ��:8|{����6f�hiY�A31l�{���?���� ?k׮�%'/��I�z� ^����Gڱ��u��m䈑2����*ZQ��oo���1�[~s��t��ǊV��'o7n��~��3�����y���2��T�	���͊y��@[�YyĈQAk��1���m����l�.x���?n��|8���+���G��s�v( �N�\i&�̩h�������J́h��ڿX����oP�>p����}�M�J}�j��68��?8B���l��#l��)�8WI���~���^��j�*}��*6�Z!����*3�~�}�����FG|�Z���v(�'s�>Z�������Hኈv��?��54	�u��:M��0�9�>��M7�\��nji��"�PKs|�:���5�Z�r�.M��N՛���v�ͯ-n��i�׹�>��Ū�`�<Z~T�������¯1�Xd��L�<�:X�Ǔ ����|��*�i\Q�\�Yӿ��X����[�j��|ǻ����"�n�}4���Y�q�i\�q�"��=�v��{�/'2-g9�%����_��3��P �پpY>�^�O"�r�?��(e��z��W(��������4��e�]�N��%�AkI�$y��m����j���T8�c>R�:�����#+�]����5O��g�!�p���1�69�o��6�l�-vک�E4	YE�fqT~b�c��~�ni�`o8����L�8�������=c�\s� M	� Ȁ�;𠾾��4'D�~��2]I��\ ��nmmWnL�� :]�a���@������T�����u�O�Zm�-Zd�������C˗�9"׮Y��R��+�܈m�wٮ��rvW�*��|�C����Rĭ(Q�D����וS�r�~{����/儨F�����A��;v��a�4�<�H�CC}��o����K�)h*��E�L�D���/�ͺ�;xr��ԁ Q����"r7mv���	���ΞZ�Ɩy?���ARZ8�����[�#�>l˖������Z	���m����Һ$}޶����t�5���ҕ�۾m�=�b�<f�� 0M�pP�Y������C˗?��&i۴e�3��g��X�D�vuw�=w��l���O�|\�!#�x}�E��e!p�e���<��@�� C�{�����:푧׬U>Pi^���f�E��D"h���9g���8<vY��G�2��:e�p�N�P_��("0r�wyp�H:�j����Q#G����\y����u
�ټy�͘6U��%�c1�@�E��������u���ѣ��M𯭉�͒�w���ڛ--�mܸ��!h�B���\2oh�yn��S�#�%� ���U~Y���Ǯ^�ڦ�;��-��ϡ�<��e�k��e�3�`�H��
��_�򾮀۾�_~M�+EU�/�V�l�ٞ���F�2��L���q![���J���$�Sy�&���f�bI�� �D�^�{,��n�{
�)>�|��`��+A��؟��a7�懙R��9җ]���m�[t�������1�������C�"rV\t��ǸO�9ݾ��/��OR6�js}�6k�4;�%���qw�o~e��P6r�j�u!7��Yv��9�[����־�����X234�U:�m��I�ޫ?�ۿ��=wڝ���n�J�s��ۑ3����':|��=�h���o��G[C�P�Z��z�o���{�L;F���_ڭ7�d3��#F���$8h�{�l��ʷ�f�NU:�Ͼ���l޼#��]m�l��f{���L�����w�}��l����D���l�ԉ��kB�WLW'{�|��?�8F}�o��ժ磌�2D����~��_��������ͤm���v���(r�r���ڵ���� j�GJJև).����*��N�?��>�����Xxc�*dm�����uv!���G��߳�O9�F�/�L��^��5�5W_e5���|��ؿ��'��γa�]��z�wi�T&�c���p��y���_تGW،#�i�������w�ǆ����c'��ǿ�����2a�d�?L��H?����^��ڧV����>ᤠ}��j�O;�����
�<�}z���_��-9q��Ż���;��Ϻ�������ۏ~�C{�6s�Z�P���X����Û�1{��5���l���,|41��e����>��?��@�����/|�V�w�͞��[�kd���W���
9f�{���\eg�y��^p����̙�>��ٳ��j��׿aO<���;f��x���j�c�{��DfLm����'W�q�ۼN����P|o}��� �3�<m_�����.Y*�!�v���/�A�k�N�������_�9!���k������m�gB�S+W��~�c{x�}�p�)-��D���� �u�/��	{����	g.�9���ec�6�E^j3�(z���b����أ���L�W���~�ˏkM�
��u���{߳�ۖ,;G�-�0�\p�M�2M� ��}��U+g�>:'�i������,�`�rv�2oZ<��h��2��|�&���^���7XM�
�^]�b-g��+��}�˟=����܁I�|�`��y]�����-E�"D��}Pp$9B���X<q+�R��?�w�z9�_)XI������[��,?Pq��4��hs�����=r0���?�/uJ]կ���?��O�95l�#+�,sh�0E��ǅ6��N�O��&EP"�a��Q#��}��iŞ6�w����_�p�mX������>������!í�o�w�����T�O�����&�XF?��Oe�1���f��x�	������?�vE�Y����!C���͙7����?�i�k��?Pk�T�<RQo��c����Z����ŭہ/�"�4.�f��0��tuC!�7���A�G��a&�m��
[����|�/��.�=��4J[TQ4XG:�2t�7�Omf��j��uYUc����Z;�A����m�I��L�!��Z^���`����&I�"`���.o밡C4N���y�I'��?�y۽�5h�|�k�j,�L���9�Erb��y�˖@D����۪||���|�6�A�/��A�V������N����9��18n��:1�Rc"F��j;f�"�η�[|�������/#�����F�u��ߛ�E(c�T�M�b��:�����n�G����<kau#�壉'��[X̎�� ����LU�U���e��_:}������22����7�q�M�v� s�2?�|545I��;�$�l���ݭ{����%-�*U^'��5L�
�W�h��w��h¹�{�����ȁ�Z[x�!�&U�Zk�29�-�ϧ�f�RO����A>�ǌ��o"���e���Dʴ����){�ٚ'��̍?���v͙������p�'�y�����F�� n�ږN�轉��6NĞ��(�s�>��y�n�.��0p{�Kqо�E<����︫&*��F��pMD���b �r1k�R�`� �Y.@!�ai/2��yP�ڈ����@�J��-AW��`����4�n����rI
�`�S�L�"��+u�'@�b��5]��T���P�R>g�=���$�r��S���QJ�{r�6�x|aDL�_�V�M��{�-嬥�Y�4HP1�d:HX@A�yis{�ak>�R��d%��?W(��<�N"�(B ��-��@�!u�e�f&c�(-2_Ɩy��� ��u�hD�[�kd����c�h,-ͭ�O\b������<&�6A�t ��؊2�"�:0k��q�6�|f�j��N�iKJ3���(bs�芇$�C�jLi��klߋ3^޾g֮��X�MGx�F�ݺe������/��x֪]���u@�|֮~ʚ���TU�����^	o �=�~�mܲE�WC?b���IВ��&���WY;i����sƘc�Hŕ6n�[Zl��+�K/�2W�I�ƍ������
M�:(a  �J&S
RA��L��<�B�g9��/f��ǺRN����u���N;��[[��"�sH��m>�?��.��r�-��&�~�e �1_KDǶ<�Z��7�s��������z���ʰV}��hyZ�P�t(���4����R���m;m����� �0��(_��bM���mxFidfRƒ��P��7��"�N�ƧW[��8eJ�)%����R ��uߗ[ׯ�6���� �x1.[�	�},wl_kO�y*h�|�Δ��nH��e�c1۲�i��	<�q�YY�yN֚$��sb��Ա�H�ן6Q��r��}���c崁E��\� �~��b��^(��P����Ⱦ�a��:/�-���LJʋ2�(�{4d�Z�l�D�;��8Ŀ���@�ghv��eU�Z�����|{
%۷�犊^i{n��gv߽wG���y��%./��c��mv뭷ڮ���:%�k��5v�9�X}����  Z�=w�}� ����+V؅_��쳖�C��o���vz{z��u�6;��S%��v� ݸa�=�r��X
r��轗��r�1Z[w��w������ۏ�@n���O���H�g�ك�?(Q�� \�����JՓr��oW>m|���6�|=f�u��!д޿{�w�\��4���.����mI$;mwk��X���������
.���I'�$g�Ν���9X���>��EF�Ǽ_��r�U8����`v�uؽ��c=���@�5#�s�ғ���lm�ٺm�=�������˔��7�sK��|.Y]]v�׷i�&K��S�Gm����,9j�"<;w���sA�����q��%	��SN=MZ��}O��Ҳ����>j#G�� ^��:�=c����ֳ�U������f��7�C���؅2�m�.�6�eo���������Ӟ^��N��N�2Y똽�}�vq�}�w�E!!�8�1��;�6�)jj��h]��G>,`K��=�o���%�w�_����X}M��|�6ml��>}��3$Uokm�'�|���_�������ź6t��x=�$��o޴Y&޺���gm�2`�ڸ��c�Ne �R>���OZl�}z�:;�9Ҏw��j����������U/>���f��B��ָ��x���f����OH�J���k���	�4��#r޴��!(��?��Ta5�w�z�Iq�M�4��c�֋��^>���{�]i�v���o��:��$�����>�i=�_]�/jC������Y>�ט���̧�U�/�l��m�'M���5���j�|�����¨���Y[[c��N�u�q�q�	e�=I�c(��{��y�בЬ�Ǚ|8������u���@�]]rh&�	���w&H$|h�*�D�U-�ԁ��\��~%6�{Ĥ��!�s��.��n��ɖ��%,�c�;ζ�p�G�m�����e&��#�v��GΗ���t��QJ)����z��e?���yGk'L�޾n4�,�9�Bidr}y�T78(����GZUe����$�C��a>g��7�:9q�=a�9Fuΐ��ر�/��,�*��;��{;g���j�F�����9��}���>%+����-��������3ϑ��A�T�Jc6z�x���K}�C�h&m��u�͚5Si� �p�/\��SɁK�⥧H(56q��/M���s\�{
Q��Z;����u��ӗ�@�<�N\|��S�zsj�	ǟ��z�LH��P�N�1�P�`��l�Ir��I�����(r���Sf��:O���FhO9m��:��CL��'Ͱ\o�ƣR�fKvɤ�cU5u���Ӽ�7�/:I�#R��-8�x���~��0 o���v$���u�堠y�;�e6m�t>b���d�`LИ���;��}g�9�����
a�>����F�/�,�	\`(�'L��;Qf߾Ȕ~��g�Tn��Z���������`��|��ψz$+F��i��i�P7T �����OTO?��u���E6��y����]� F�gg�{��?�_j��:���jr�F0OeU��w�)Km��) -@ҿ����s��m�[�	�K�@`�5�H�n7o�bc|n�3�fΞcͣ����z[w[Um�]r��&a`}���6hyv����.x�uut-������:ʚ|��J@θ	��W^��+��;k�^�VQwd��B�a?sꚆآ+�`Xw�u
�ޑ>O���ZF�q@�*�P�6^�>����a2�K�ҷ^���F�������o��I:[ �&����,z.g\,gΚk��-bb�/��7���w?G1�<��X"����ĕ���i_��r��K�v����0p{� �D5���_H
�ῂ�Qi����JL��,�t�J�9�'�V�A�!3{�ȧb.h��r�t�Ne�68��m�=��f���(@���W��)�s�t�'Np!4U��ȸ��`�s`#_��:�W�9�X�l�Wr^j�vY%�N˔q�Bsf	���.q��=ڏ�vO>ks��uau�Y���B�0D�@��sѢŶ�������@;��y�����w�|��D*!M@�����ڟ%ʢŋ������������p谡����@n� mZ��	��e�(Q��.�E��Ш��K�1�uvu����YG��O��^�:HwTK>��t�Y.���>.��/P�e��Z�.%AOUD�?�7uƴ@qP���8�D�@@J���9 ����&o_O��2	W;H�2u�4\ԅ)a���_i��M�cO{�L�aSf��x�@�Q���g5���3g�9�W8�cc. �hv��ǌ�7]|�P�" ���@�V�	��XJh0i?��n_#��.4��b��2}�_N�kMt@NW�9AѲaNO�; ���`�?J<N{ҩ�4�P� 6� ��ǅu�/Q���\0ף=���*@�gh��k3����C�6{���9-�@[غs��'����u'O�؊@~�H���?�t��ǎq5�Bee��KW0�:��}����S��hg.;[�����:���,��q9���w��=r��z�B�V� �x���5b�H{�[��zGC�4E>/�Ȍ)�]�Q��*c
뼂�*�<���L�r�8d|-�z��ڿ��"�C�_�/��U��[��§��"m��i����ܑ���뱔�-�WD�a��:/�'(QL�"-��A凌�9s����(Ц'z�#ߖ��x\���8"t�4n{|ۂ:Yi����t�	�r�" ��7 -�!�
ʂDL  iMD/��v��GĚ��D��C��  >`�爊� Ј���y�L���0��|eFX��v��m�LC}�t�q�̃ G0����"#Z��C���.��U�iܺ��J���f �P'�$���. �Պt�M����n3�bZ	�@��J� ��>HG�#�K�_>� �x�O-
}@k�_��a�2Q!�ksh�&%P�X`�Fx��%�҂�����˛�ƩVs��c����� ��U�\	Ի�G
Ek O�@6[Ap.�@4_�FMw%��� ��oL��7/�4 ۷lV6@kz�	hp�b"��*ѧhR h���ȭ�c�'�� ��FAÈ��N[ -�����E��h�x/ �5HݘS{���_����u��`��=�f�R!ub@�SѸ �Rߤ�Bأ�G��B#U� ����ʹ��\Ba�&��L!�N�Q"��:�`�e�ڱM�/�	�����P:���'G��>=���@o��#D^W�}E��X�I�V8-d�X��ſ�q�z�W�Z��~���w��e-:��h�
�M�X0�v���@��E�}��WF�Z�J���?�+֤�^�b�^`ND��m4vw�i�k���p�	��8�����7k��7p����a��:/���R���	�J*�����%=�T��:�}\�K9�=Q�Կ�VRo"+��. �-A�ƍ!�-�¿�euA �[9WD2����O�)7rqIt\pe*�Bz�R�7 �C�H���B�"t9��ѣ� ��N�G�e@YVa���M���>RP��}@ے�����וD��  �{0sB��eh$(c!Y���@��%
�4�h@� ��-B�͟ï�EH?mG�ӶxE\��',���#�xT6�GZ���%��z��}@�cj���1G��|ԇ��Fi��<]�\�~� ����?m ��ֈg�(���"pr ��� ^�����R�ۛ�\
����^����u�١^�(����������ؗr�XT�ցI�:) �x�o�T&���~�R|il�)i�XWU"xޡˁE��b�A r�'�m�:��/�i��Bi{G��T��-��͸�v��T��`��|��'*5]����! �2`�v0��`�/�����q<��p	j:L��4!Y�I#�#@ѯ��9��*4'8����a�<q)! &) F�R��� t}~�O�/��(ptق^PU,�te_��#� [K#J��NWg��{����5��o4� _�T�k�k��:S���1�:���.#�9�K
6Pƻ��6�m��Z���{���������B�e�(��C&�s25@e�3�������}�*���^s�P�n2�k��'n��(DR8���6��F�`�:�t?g�����`��pp��.�}ѷP_��V=@QG\q��4>h�H	ǰ$��	7��򟱒�TW�&m��/Q��SV��_�Х����)LP��](��~��GL��W�R)�·(�ȁL�tH��Je����f{�%%�9��PE�D"���	��e-\e�Z���/�$L��I�@B`��I.�l�a��R@EZ&
�l�����2�Kә 0�c�+�WeU��)���|����w�4�d|y3 �~2^e�+ҩ*�[_6���2K`�e� ��	�2/�)�Ja-8D`��2%���ەˆ(a�P��v��+'���<љ�U����򥠡�w��.#�8��L��S��R0����BS�`�!ؙG��?6Ɩ� r1��*��|���`��A���uJ{���5��{���G�}�6���L6h� j�����b�����N�v����?K:%4`29���Bm.�����=�)�ץ�`Kg�@?˸����W�s�u`g�h���E�W }������W̀#L���u+�����o�\X�a\��n���+q���g3E%�7����,���w���8�ܖ/l}��+X��!]������b�_�4��t:�0�\����b=�{C2��rN���C�/��e\L�y�Qd](z�Ѱ����;���*�s�L>7�^��O]��t\���xA�d%�N���[m/W��Y�K
�z)xĈȤ�H���P��+Y��������|^��)S8��^��*�4y�p)Tڰo���폩�2F
��Y��#�������i{�J ��H���4x!���W�����Bg���{�`�����ǧMc	�'>ThN0�aF�@������ł��Z��(� H Iz�e(�`���#�&S�%T�w��c|Ɓ,��!��f3k�����PBA�!0-�g�` �{}}�u�P�����a_��6�z���٠=��$�Z���=G>G�e�����
 i��Z�^G 3/m�# ��K4C 1�DR&�`z�w$��!�!�ZU�>O�S���ɼ��d��	��z��䡉c��<a����+}�zL�2kŒ��g�k2�*
ӑ�`8��&@��3#�cż7by�h6�Cr)ڂO��}��V8��E�i��a��Ü�-�fLi�x'��[�6 P�9�ː�O�=&l�=&c@\t��!+���78�Yg�#��@@� ��@i��%+�N�f_�����5�~���_3̺�/�8%��
�r1ⶋGր�+��׉o"�����O�ha
EeƠ�d,D��d����-ej�q���YtH��a�P®\oWwgȎ���4�\Fc���O��}��PW,�O����Ƽ�|s��m���]��5^�0,��w|>Y��ҕǠ�����*߲��Y4 ��aV���圡�Lk1�c+D>�2�s�iq�Ͼ��Rl��т�_�ܼe�l8�G���a�v��HeU�q)r|�[<@����8����F���j���(���ԾM��0�ܚ��!σ�vi�����Z�},�Ҟ1I2B���%�l8tᎂ��eE�j@S��8�;Gt 0>l�8XՓ1�44O:��Y	l�Y�E���Ly%�8����->T$�����\�N�f+�q��j3��@W�����>�u����kQ������8:�I�M�(�<�� #�& n������-�8ih��A�R[S-�A���$)��ǡ?V�D"` ��< 	aM8��K>Gq˹����Ѵ1ƌ s.�.9 @#lh��S�1��0i{?��BU��D�xm��� �r֙��h+�j	4E9�?���9#lcֹ�#�+��Ax*�%���+��^H}� T4�8�"�,�_uCm��x;h���YWר5� LоR);|�W�)ڬ��d���8_��JZ23LƳD11�q`$���wf\qZ	�E�mk͙d��V4\ M�� �tL����=a�
Iu̬	���k������S�6��;�����`�s.�� ^øL�s/Z�b.��Z4=�	���
�DQ�s�Hj�w-|��/�%?A�K<ǚg-) ��U)���J��hU�]E���%��*�y`�s��ҁ��|v�o��p~�\��E�2��1��-�|ڨ�/���"���T�"NF�bȈC����W#Wi<;��F)����#x&��v���r���h��>'�v�;�HTʤ)���P
���/���p�)��/T���dM��u�,�G��|�Z��X�������l��+�B`��2��(e-�"C!?�F%8�R# N���8c;�PX}<E��*ϤR�`ZL��O�
��H	vv���LD$�g8#8`>IT�t�c�`-k�dVa���8�Iֺ�5h���$3Jz]n?<�P��䛗��S��L��~2ɚ`�!�����_ �C 3�6i]�sS��b�`��"rK��)'l�g�Q�pNd#��I���b���L��B0��ʁ%A�0漽�� !!M_EJ;�	�c.�0�#�PT�u��"?Ŋ ��hN����*�S ��,�c	As__>$@�L��nA����0�6-�^e0�z�К��qÞ�>hi�?ڃ&)#��P�G9�Ѐ�H�`lUE~�0q��@I�{u9H���x0!�X����#�����>%�]�@�p�{|,zh�8Pd��T��a�E���E�ʹ��oe�hƃ&ࡔ^��s��emQ!����ˊ
�� ��/��c�Ǎ}�3�J@>T#��r��"�8DE�5>�x��d\e=��a+�i*d�\����J\�CQ�:�TLu��#x�ai�SD�wj���(�``��1�	V�FZeL���q�2.5y����i)h�������.��/^<h������N�Xd���a6�
�����g��nY^,h;X��/��'���C.�9�̚�2�z�E$��@b+z?�����ns�y���ŕKp��".d��{��z)�C��uO_�_B�B�C�­��*����@��_�ơ��u�fkl,���Ь|�W`��7��/F�C�� ��@~:����ln���{5^!34T%��!�-!̈́��b.ȸ�'a�s�H�����I>P%	*E�F>Q ,����e���UMJ#H:�I�%K�(�]H�Z>$5�:�	�	ZR.I��������z	 "�$�P�����#���X*�:[Y�C^�Z������b�cLäü��U����^�R�>o�]	Ҁ�0
���@��sa͛�:�#��;�>wh����O"k�qh�� s*�%��J)!�fL�5�E]c�.����ֆ����$�*��
�2�ge�H�˃"T�޼���I��X�J�L�̢�0΀���F	z�p�&6눴�� (}��A�=�����(v�z�.�SV�|�'y�MX^��@���}�*�;u��;����Ct��E�1x�zq�=P�����������Y\k6S2M�~��׸k�����ځ��D�T|R,�<�4o�Z������H?���2���V�y\#���>j�)^.'��ơì?K*�w��{�z�M�������p��I�sH���`��v)C�)�F�ih���)�s���|���p�̣��2bʰ���S�v�Ƥ�!M�� �1�ա|�e��������ʠ���{���g�8���R��
5I^@n�1i��R���D�["�9��CT$�+��^B�����Ó��w<_(��D���<Fhz]������=��W���s�1Gϗ����?s ���t��S�}��48�r�?��i۵{�L�ޮ^[r���LP�ܚ{�e'���V�cF��Y��� ��t�n{r�c�c������6{�����:!��kV���S�k���i�.:���u[�}�����$�)@����yG���D�ѾUO>����l��!��_�5u�<m˦Ͷ�e���{zz�=5j�͘9K�
�	8EK�b�r�+ ���۾}���~���	�����>f-^'Z�wcS�M�6S���� q�soy�6mj����:o�� ��w�� b����V�s��B�)Ӧڐ!�e����Q$�5O���5�7� �q1r��D ��>�����|n13O�8I��+�,d�صk�mڼI�s eÇ5��� �=�j�u�\��u0r�(3f��,Gm��	�#�%�Kv��ǎ+_K�����dѲ�Y�	21 *�5;ԁu1'h-�;�m�6ev��u��O/mUUF} ��5@k{��1�s@��Q����y�}����co �F�3cǍ׺��p��ӏh��*x�$�4}��<2d������{����[��)k��M�:��Ѭ��$}نg�)]~d��'��#�ڸ	��(������k��R�IS��}h�p��uP��c[�����C��Ys�yD��w�[��M�y�f]�+�T&O�b&N���ں[����^��u�����P�g���[��
�@���/�	S���f��m>Ƥ����1��7����Kk��J9r�3cɺ������qۻ�;�_y� �0p{�����@�����`ɮ����A0����l�C�M��3U'uG)�U�`HT����$CA��-��#`����V�Z �5DB�7�篁0��{���w��]fLUWR�qa��)�m�{�����&�a����M�1S��Ѳq���{��n�5$�����M:�r7muA ����~�[=&4U�]P�<�앩 �o��o��_߬��E�	��a���7��'� �ܨY������25��_����N�`��i��0�P� ��n���7�!<b�(d�]p���\~��EP��v�M�P:&L��� \$���F� 
&�;V�nw�njiX��E�'��h��V��ֱ����g���o[�!S�N�\oN��Q"׺ ��}S�����k���z�l��bn��Wv�����c��%՗��GQ������_�֭[mĈ
� Zk���!��6$��\i?����>\B�����ox�4QP� :�|�q����'@�uJ�XB�����ێ�֬zҮ��;��&MHa,�xە
\@S��h��������h��K��R}�C�l�;;֬Ze?��g.ܷ�x�c
��_bn�h<��u����vV�O�gٙg٢N��6��a�쁻�_����2�h��65�$���<��c��[n�g�yZ��;��&���?���t1b.r�N�8 (��\��s��S!Z��-��7m�(�/c���|�R���}�����~�˛�Ҳ��md�۔��#o,ZЕ�?j?���� X
m_��S��+.lO�|����Nc�&�^
�/J�k}��c�}������K�3��Ș}?ᶲkG����Sk��n��?"����%�^����^YUiO?��~����꧞�)~���B��{å��,{���ۊG�����W���E~����X��qѶ�"�'E.�^y�6p�/�q��c�l���l/E�y����r/��A�8 me�W�^�;��!�?zϠ����a��MM�?�b�/
���/�vD����s0��#����������@I��v�ú��MfCn���{�}���؟�s0��E	Ϲ�b���Y�� ��믷��=�N=�,�����8�7����Q��k���.��r��˴�`E�0v47����u��E�^j�\v�@�I����l$:���o�{��ڎ;n�L��YqЗ��4��>�¾����{��;���T ����w@B����_��|��x�� �S.�����X����v��Ev�Wȿ ����
,J����ٛο����H�^Ю�)I��O���,[v���t�R�������}�;���@�i��a�Օ
 � o������?�����$;y�)V�@!p�e�o~n�ɟ���}�N=����|Ts�Ta�(����;�~�[�p��y���2(@����z�9�/|�?}\��/�ā]�4Z�s>h?�M���^N8�D;��3-�뎔k�>Pz�5�6�S��;���#��𕉟)e�1�o~뛶p���?���G����s�����+_������	���ތ[m��V�xP��tJWG�� @�w��:H��׾�\�W_�~�%�� �5��eC���g?���&�;��.k�}�&��2� K�m��W���	�W��F��y�.�z�헮
�����}=ϝ;��󾫔h H��=�<�v���������\eC��پ��9cI�:z�����_)ˮ���ڨ�c�ņ�LgK1���f�Bq�%�X��p\�¾何�5��}�??o'M��������1lP���)�:�<������7�1c�*�I�����z�_&�;����7�z��W�%r��@�Q#~��6�]���$=`&�����a��X^�Y�C�n;`۟��̅��iK$$�/�!�����*�������~����O���6���"�p��&ʛ����������c�g���\ ��k�����\ E��O�f�h,�Q������{Ʒ���-v���٬�3,��0!�2Q[ $LR���~�ܣ��II����EE�@�8�oj�h�5���Ĳ�]�ceMƺ��V	����o���e�����ioGk����H'eV�Q���-&N�da�B(uە��q�#��b,<�x;i�R���,�P�����g��%��	�/ ��K��L��s�!^_Wi���&�{�|���OZw�#���&�S���l��( I����hG|ܗ?��u��v���!�`��mhj=��e�i4/Y"��ˁ�Lj,�8��~(D��6��ٶ䤥��G0	��z׬z��A���}�X,�$)���{��������3m��%2�c���������B"��۸I��s�x� K��]�Lu�r����?�}w�c'N�����R��UH����?��#�����>c�vl߮�uIoV� ?�1�;�S_>�Md�w`�ՙ��k�yۻ�}�ɿ�1�÷��Z디aDC߿�^�0f�?w�5�����;�ց;�#���"#_+ ٺu������s?2w�3L�7oX9�#��h0:Ȉ��k����e���>d�C�����-���<ZI��7��@��i��?6. �;|�h'�Ab�3�-�S�sM.&�*����:����:|,N������M��1d}�|��غ��~Μ� zܸ���>�LN}b,�x�qif�x�[v��;�C)��iԠ�ٸi=n�v���z�22�wv��_�B.%���ز�����'��F�n���\����ɒڸ���q�ҥ6��l����,M$Is��&�_S����?8hؔy%��xS�rb�}�V#�����9��:���!׊Q�-%Ej�����j+ǖ�O��JPL.R���ׄ�Ky�MFA;���x��\V���ۯr�/!�^��z�`-U���@ �Ͽ˥�yؕC*���ͮ��L���G����6�s���Tz�8��r�ߪ�V9�9V~\8��);�s(D�����UoM.���V��� �FӰa!�����Ə;�p���[=��� �C�y�����ڎ��)*���	h�rM�]ؼi�M�4Y}mI� P^4��-����s%�d2��jmk�Y`E���� ����9E'6� ǌ���- ! �m�w58 0u)XB�U�� ���ϭX����]8`~�;L	�O�/<�v!D�{"@�x��Bp�w@K߰��!�i?��mQ��CBw�<�vn�&��s��%��"A\2DD���|DD��!�i]S"�����9�������3'�<�y�ƿ����O�K_���L'N�,[���C��Jq�U(��V��ii�
5	��c��ژap���#�؀�+%Wg�٣�����k'���J����Q��h��F��� ]&Ȯ�q)?�������`��-����Y9�6!�pA��vݺq�F� �.@J@�7\Wj�w�=JQ��އ-�G�L�'W�:]��ku��������0�Bą&��ݭ���y���œ"�~.�6XÚ�k��/x�wǌ�=���#��`��	�蜅�D������3���h�#��L)�H�5Fn\4ω��o�%��	`_\ ��E�.�W�U���4���� ���w�Ԗ1b�sv���`���u˾S�{�~�2��_�?��(�40|1尩�C�)!^@6����-�i�� ������O�u0`��n �����Ge1x+Œr!�X�Cdg��X�p�mbp)��z�sl�-:<9���w�P�"-�H��\��J��G��ڀ�{v�;�Aǘ�cux�V�Ŕ�m�eKK�L@[��ψK-6 �x�c�=.�8� �|��rف�Ku.V�zRz��1zJ�AU��۱m�|��L���y\����8NQ�(�
O�T?��Ў�3�����7�G���8F�AB l��(�B^��j���>�@�B�5����]\h��Y�
`"��n���+W:�lU�w��) >�E�V��h�g�F�{ƹE(�,  �_U����!�������ත[�хmE&%m�8����h�#�zd���F���v�ۥ�C����w�5��.Z�?+-�-%����X_�D��-��x���y[��Z���qܾm��xI��e5�X�V7�7ꂲm��>s��=�6T�%���Ҧ���ٰ?"�<X � kL���Pi�%��6o٬�Z1�Oк��(M&O��q�5� ��s�!��|>�z��B�Tt cp,�Ce��#}?�j�M�4UQ<q�%�1a��gLgT�vz�8��-Q-��ٰa���ki��jgd��]�ъٛ.�@�/E�EE�wiN8o�Ƅ�+��#�: n�~������`Q�D�(�_mO��B���^1:��5a��� =k��P7�~W�͟�����A��3V>˗��y�Hې�y�ˎ���4$� �?(��?���@�=S�[����W��H�F��
�@��zm�vl��:�f~�s�H�Qz�i��`�v.�`xF��t�38�|B�wl�6��Ri���� J��4����g<ϡ>j�h��;߱?�8��#=S�Bi��!z!�(��}���������Ƴu��}n�h�$d��;����O���4	g�y��e|�9 �<��� ����������=�<8�zo9�O*"{%!9�ޟ������Η9�Y��p������[����b��ԧ��O��!M2[��Q� �K�����o����r� )�ӭ��I�2v�8��Ol_��m�mD�i�v��f�Ǐ�}�6u����?�	;��79pjphua:l�0+��|� ԟ���NR$$`�1D�d�U9M�̞����0��:��]�zIw'�$$��0��:>A�������	`FA\X����̧�7�e`Dd�O�|O�=�e�u�,aI������{����Su�֭:U}�RU�����tW�{�g����t=]|��0@��"�#���}�Ŧ�O_����S�{W����ΟK)+�m���X��֛�,�y.dН��x�C����Iz�!���:���� ,1v`k�k&F��~�!}�3���x��mk �#ҝi~w���V�j��BnV<vp3��ⰰ3E�����s�A84@-��:�h���@�|��t�����fb�Ft3>�O 68���@��{��<A����[ �;︃�{ᅴl�2��ǧ�r[8���
�?�q���_]��t�ʃ�u�t#6�h[���v}ﻏ�ݟ�,�{�y�6�q�� {��?p?�p���m<NaW9:6F�:nK���}���._/ �R�Y����1��;�^{-]������(� ����>}']y�U\|�1ͪ��1L2<=�����J�o8�����{A '�uњ5o�q]|�%����� ��j��o��6o�������	��!��m{H��k?�q_,�cdl�%�!��"�܆�/��n���ЈX� Zp����"�MJz����о� ��cVaMġ�Q�jUn������g8<n��q�~K����A+c�f�mU��T�P�[1Xz���:��=Zzo�	V�	9 �x[�e�މ<;Bl{q�+��f�idr.� Z!�-ޖ�T�Ė�bK[�Kg�`97v8?j�9�h��a�e�@]v�����}�z�fh�@�y�-�V�X��z�������_��=;�rYs�Z:��ch�ڣ��X��>��������O�G�?:8ȱ�n��&^��AEz��g����~����\ �����t����dx#>Gl�0`��G���y~�E�A\�a3|�������M������-_N��~PC���w�_��:������G�|�z�7�b�<��:� ���Q4���3�`���?�1�� Q6*\���<oP���o~��l�"6f? �ǆ1������������jp�k�G6\� m0u�)�ҷ��W�e�f�K`0�d���秊�q��azʩ��w~�>��h��^� F�|�^'�'�+���䷊v��oӭ7m�M@	��e�].���^x���5�. ����o�cn���_�:����ǟ��	x��7�I����<_��-;`�~��B���d��q�����6\�QZ�����?�mm��	��@���W�B�}�f�`s����\N�/�߷q+4��#=L��8Z�|	3i{���W����[�@���`q�}�������!�@�|�{�Z�@@��sΥ�?���Pp��W�߁��t�G72pǜÁ��G?�!]wí�h^'͟�O;vl�~[y���^e/�Dy|�~y�E�(�<��vH���7���'��'Dy���l�٦s�=�^w��x����N:���w��@m�P6��j������u��v{�n���\���\��:�y�%fq֝t���7r�[���SO��X}���� F�t����q~�m��$���f��bw��F!�� �w����� �W^��]�zza�</O8�D������e��'C�C��5��H`%�\������}b��=h����vXG+^Ɍبh��O?M �t�M��|�?W��B�&P��8��#��*9�J�'���C!�e��Q�9B�>�`*x��\�r]�0�*ï�~yv� kl�E�0�����Y#S=�tڠMEZ�tC����Ќn�pynh���98Y�W���Y�t�;YzZ�6(����F���P�"��%@X� "�����A��>N��J�+���A"��i��6�(羺�3+OZ�j�Bfh� I���X�o,,�0h_�d)3oP�����N�5G������o�!��-N�lS#` ���c%���KEUl�����M�6�믻Q<w�� �����6\U@����Gh����i�#,�`� �����1G����	���D<*�@��������\O;8u��@\��*FD�,_5�j��t��	 8ĩ�������ў=�m����b��C���af�2�
1�8;EO���<~�������G���9hs�~�(�
Hs��A=������vwҡ���֯���w��  0h#|�|�_?0L�{� `����0�y�MX�w���(;:���ཱ��8,I����Z��>y��ܿv&p�Y��%bSʻ�U�]N;�%� �P��b0����!Pn �`�`c T�� ���p���.�s�;�^z�Ej`����Z ��k���p�2�u9���C��c��{���������L�O��Y�6I�7�r�E�����[10Q+D;C��� ��{��r�K�Fd�� ���Ab|R��[���k�Q�7��2��0��N<�Df/sA깅�R���D}/��"fr�t�y��q������p(X%�+��nhxX̙������8sv�8Ty�h�}�_ �p�� ��7��\�qo<����� �̍����L {�{�y����k����h�8�p�ML��w>{,�q	{x�����M���O��CW�i�`/����@9���S��-<lF֒�2�G�=�BL��� XA�{�������,l;
G��1�a|e`�A�/��3�X�#C"j�� MC�Ʀ�q�W�;R3����$�N;.��wN+ ���b��\�D�����/�����_����A�3�/���򡿣f����'�y�vT.P�n1��(6C��h�*��xF���	�����z������.ۯ�:C��8�0!��iv�� mϿ̮��!���,��h��������Y}��1��Ɏ�;
FȰ��I*��X���7�ΠJAܩ^�홤C9�7<,�0��Nu3��g�����W�w� �&�-BB@݈xl�ă�?l��hb��F#��C�L�|�I��	u���L�2Q��y�~���;��O�;��f�g�^Z"�M�Mqb�<��"�ړ���'H��<������r�ؤ����{�ƃ��-V/[M�����	�&U�9�)��*-  S�"��q�P�;��NNP������}ɛ� +>��_4Z?l~pb�#���T�B=���f	p�d�e<^п��<h�������t溸]�y���1��e�K�̆��*� � "`�m�����=c��F_8��q��;�~(f��������`� YW�b��p|A8@��phg��^�1�\��{��|���r�["�39{G�p9@! 'r�!5�4��w���0+�}���1��Ę�g(�c��#|�x1��y$��;>taދ�r�>�s���-�m�ļ���&�s����f�%B���!�i�|3��Z��c��:r&3�������K�`�&a]���9�;c��+�0���gPK5��/,��L�c��g<�ZrMĸ�D9�t��¶m�Զ���;-]��%�:S~�h=���\�K�] ���ς>ā�s�Y�&�G ��!�f<pS�z<ht%�m�"��@p��2`�[AOHל9|Z�Ju�SϾ�!J����qNB���{�N������'���z����a$�TS�^���)�s��2`��z�� �`Fe=����ɋg�	R+��b�ͷ-.�_���^a���g�iؤ�����=�o߱��#3e10@�\
*<�%���k,��/<���}�u�{��F�ˬ6�yb�~���NP}��� ��\���K��aH����Z����%�ϗ'm<��j���`�Cp��!7���&�B�4J�hR��A�x�?�අ��16D����@�o.Y��  �e;(
۾I?^�6	�
玝��S{D�`���k�|���XU����;C<�̳|�d6�@���'�`�U��� �%���#���~�ܠ�~،������d@�9��(������x/8s�6�{����*z�c������s�]�8B{������<?��=�� Gy���.�#m��'Z��ǵ�����;��`s��Ęz��f��/�gт~f�8�.�j�1��w�<��AV��~��>�� �},�[�U�*���1�����@ζ��І{�>�m�s]|��Un��uC��~��w�$�c�k��W�N��tdM����[C⠆w���D�q&
�ѩ�PB��3\�ǧ�fU��W^�w�Ƣh{�L/l{��:�Nx/��W2�8y�Ϭ����('�p=D��y��\��na�Y<��f@X���SO��ݧ�^Gd8�Y�r�r;�����y>����0p!�4���*�V�q4�����X&��2�a�NB5���T�ӧ��f:j��r"��B�d�O,8�x�88-�8M�b\u�A�����	�E��F�w�����#��d�bB ���۞��L.20���lឌ#�U=�˭��O"�$�H"���Y���膮��؛����[�<��F��IV��ŗvq*<�v� ^S	���x�f���Zl?�
�J3Q�N����g�A~�u�f`�N�tX-��g�y��d��¤ p�Ę���p>DM��Y�����&��Sn2��=D�� ��f�
����ث�S7�N��d�D�&RI���=�"�:�ةxM�{��N�f`o#?��;A�+e������'n�r!ՀÕfCeY����>�e��s�b6y���.?��G����8����-C����R�]p��aFJGz��H\]���r�Z�{�u�x�W\xe��m��W2%x��p��wyP�L_%�{�}/�~vܻ�շ�w�߃r���J�}�I���8��^��%^��<�<�\µғ\���|��G2�C�}�s�Qm�r�,96���ʕ1�bָJ�qw�\�������D�7�����^�̔2����cG4�Z_�M�����!���<M��4H��-��Y�\������b12p��c�;�~���Dɮ�n�m�@��3�r%�=O���k��'�fQ���]�a�e�)���7���^�+߅���hUY�U�\�`�>��W�.�\4x4f��FƟ�w�J1�y����E4�z�^y�4�F��������$K�_[��H�] �@�/��,����?�]yyv�}�XN������޶��^���e�;�{d�{u���E��ޢZ6�B��Ș�߫Dn�2��̟p�:i�G,���%���ɃQ��½���;�8>�̸����Q%������ gm�$�aQ:<��L���#�+ǩ�y� �#s������uJ�%�p�4�mY�a5��eeX��o֡er�Ƹ�l��gL��l�����,�U���N�^>n��K�b@��	j��m\1�޿{�:��c�����`@���M�`  �Is:���k��+.�g��S�=s��!ll]O ���ƩlA�՞�DfN�$Q`!�����(v���WW����7
�
�����d%��QƃM��! �!��.�bᷨ<�C�i��^-��Z\�n2�Y�}�w��$,A�
|�R��ɲ�w��0�(���Z�`�书����9���&\ʍՎ���R�Z�g��ǁ��r�Y�e�H����h��T��"qs��rK�bF ���@�U ���3|�:]x�����Q\���cKes�?u��A��`q���"�-�l�oQ�6���A�K�Z��p�pP����d]Y��hZ�v�f0����}�}T���l����$�ͮ�N�@�K��?���{�{��=N��QfŦ�q�@MN/��j�z�y�Ww��^{����r~E}'�t����vC7�BPa)�>4���Q�D��cV�V������H(�$��ы�
�߇N�Q�Xh�gI���|~8u�딦��bc�DٺBUButB��zF�Uɽ1�sB�{3!�)�-�O���W�Xa�핲nQ�)��s��j�u�����2������ni��Q�1�W
,���Z�Wk��ϊ�����xe�-P5	G�c�0Or����Bf	�� 
ׯ���p�S��k���Q������R��v���\�]N�#��qچ�zy�g���M�TךՆ*e���$�-F�����VzN>7)Nu]�B��l�����4��٦�W��q�_�]����}��찀��t�
	���\Lg�u&-�o9=���I;wl�
��+�7ȉ�-��ʌDf��-IM%%z:�K"�S-lA��B#c�Qɤ���'�pb=��0S!&M.��`|�0�q�6�%��pڱ�T*+�y���0#�K����|*1 /�ٔ�����g7;�c�z��<�/�;�w�e��5X�6����(���E�5�v��^-�~�SE�wkX���:���Ǻ�*`��y�E�q��/>��طJ��єA��sB��rF[m�%�af��u䁣��h��f˾`���S�~G�`wm$�	�2��-\f��%�
+P1����J#�CޥtW���q��.�����������6;���Ȥ�����2A��9z�O�#��џr�h IĆ� C�2NQ# ���0u�Ҝ3�AV�������DŸ��wk�[�H_D�K�6�k�]���Ҧ�����z4Z^t�D�+;�S�-�R��օ��b��FH�o��A��Z9]Q�⾫ז)\F��T2���&�c�r��M���Ė�C�[��S�ժ$���[[��J��X�l~�l]k��Uٸ�ˉ�����)���Pi�`���"kX:���U�JS�a�Zm�p_;:&LE��?�����5@��`�`ȉA��ϑFJ��tς =�P���v���~��QwW7<��h(S�v?��
/*��K�@�D��8Dj����kHQA�~�L!'"��A��cEE,�w>2���I%F�VRɣGJ�`�}����*�(P���N�!��J�T�n'_��֪3W`���7�j֒r&���^�>�uw�?(�kSZL�p
��@�_W�>Q�,�
3q���<�b�E�Fgapv)
�e9��m7�ө������1nQ�8��-��6c��T�I��<Q��T'�m����s���T6r�l<�ߑ��vzŃ#���]���ӵ��R��z�6�8�����(0e�19q����&�>q7B��<T6YG��hWA���i�DG�oC��H`�ʌ�s{?�g����gP�c@ɘ�삌��TG1�~�t3dw�P��Uq�.{~���@�'�Z��v���:~�m:RTI�ɟW�éj��Z�<��qɵ�W�Lu���S����[�[�߲��'���6[t5���<Y��˩zM�R_���ׯBX �)����B۹Έ���]��zE�u�1ձ���f-!B�^�ǶUW��9N`��P��0?0�S�CM:ՁT�
{�6b���2��a����Z�HQ���Oˉ$�H�K��\� :X���`���Op+3ll�VO�n���Uh+���m)���"@�g�>l��J�U��H"����mv�Odv�t���}b���ga�
�VK�U]�5AV.W`�R/}��Tk%iw�D��2[��[]�,S=�V�}�V�n�Ɲ�x�jF��{
�eqP���*���Z^i����]�wLe2�b<�zf5i�ť��b�}-E{�fo���h��6�^u��~�}���(&�[Hj�}������c:�j;
��<@g���&���2]�v�ho��H��L�u�O7}�aq܌6��lSa�TA���j"Le�u��A�)�2%�r1����T#Qe&�F�ϰ�'B��ܬg���N��.�f��c� }���t�ԕv����Xc�)a�I$�D�_|�ej����9ȿ�	b����b�ɇ��I�P��j=QU���L��ZKn��Tڔ�墋��Q�z�?u˨eL���k�_�m�Z�6Z�����f�<wf;�3�FM��V%3���7gg�mâ�H�q�;%p�En0���ɿ���F(]��s
�?���M|�K���q�uX�?��5�[i�5[L�H��Id�1�U�ɺ6;�Y8���u�ъ�Rǫ�G͛����H	`K$�DId��L7k���}j�>L�3��7���̞Pz�[�0N{�F��v�ZS2m���6K���/�L}�b���H���223��1��8?���t�[�;{��jm7�����J�1�٣*2n�eT�~E�	{��م�Yq����T��3X�b�Fǁk�x�n"m,�9�5����}�S��z���T���@Nxj��J��C@��|c�fk6
�MW��v3�yK$�Df���u<N���t_�o#��30�M���Ͳmr�Yf� �Puwf�*ʾ`�I$�DI$_�J�T��,2�
��(af3 ����AtU�t���tT�J�L�I��fc:4$�["������qfrP/����jc .Nj�To'vV;(~��n��Md2���Ey'O�iQ>��������˻�-79�1ݺ�{h||��t�bQ�WK7���lq�=50�jӝ���X�H�7��.������k��z�l?x�ތ�f�?��g�80kv��JRk�����)�/.߷�|>W�r���g	0	��i#-��G�.;�����r�<�);�Tv6�-�f�\����O���qpw���:�`��,��5���l�S]�uo7&N�0���MM$�V�vf�d*@"�R�~\/��J�>�ř��Z�����i�Cm�*`;�N�����0���R�3f�Z�NdP+�4Ӑ���V��0#�Yb:����	��#��$R�$s�9R��a))=�ନ����4if�9�N�h2 րs<�#����f
��m��]����tG9:2�jR'�gG�2�C�&"�J�l_3l�:�l���N?�����ǥܚΰ!Ͷ�I��%�H�d&|���i|�T�=q_���U�
����O�y.2�p�c��j�� ��M�����N��J	d�a��Z��&�'�\*mS.��U]÷��39���JeƋ��D��
�5,�`���K'j;�M�Q��D�����������4F������q���o�m��{G���:z�n���]1L������Z�q.����7��U�� ��mٔu�@���#;����7ˢtG��Ť�Y"'�/x��$�f��})�`���-*�m����<��V�j���h��z-q�1�&�L�������,�q��e W�O��-��~�x���&�L+�X+%� T�{tt�PWg'�He�yi;І�Vn�MFE۲Vc�� T�fiQ������3�DId������D�e*vkS��}F(](�H8�"�g�A�R�9�R�M�P��&�r9�w|3�ɐ�J���9�G
��( -�w��AN��E�}�$m�$�4	څ��j���H"�$����������Či��n��/�Q��(�}Q s��d&�bwvuQ�N����l���o��ϟO<P<�׵������||��mq'NG7 �̞�?�52]T����:eU��z"�$���J�h�Z}�����o6Y�So��D�G�=i��U��9���߫�͞��w�~ݏ=m��=����T��s´B}�ފ�W%'N�y:��gvtv�N�,�,�.�{)���� [gG7�g����F��0�N�҄�"��$'�SV��Qb-<��21��S\�����d�藫��3ݠ��y1��l�W��f������W���6�Ư�v���M�������&7�=U��s�|��z����g�/�6�a�����G��5��U���������d$�Z�t�JY̲Y��m�����3����A �Pf�AWڊ1n�ԙ���0��K�l�0��s��G;	7�wD��]6��
ߕ�?�)����甃C��غ�������r�����\�������E����R������ઃ�o/5uQ�ߍ�*U�?�����{�{/�|��gl�r ���+D�8ΐ����@���b"v�:�}-���:�����C��Icc�d��*��i��~���2����M��?78������U�\���c��@�c��X8�4�y�nC��k�Ӧ��*F�Ѣ?Z[բ��q��D��֢���h��U{�_Cs���h���TڔŤ�3j��
�֛�,038�A����Ryr�z�J�gB6��U��)�X� ���Y:��I�F�r��M[��tWF0�ݘ��9*�-�@ۉEsL��bS�{���ԠFM@�/�jĦ�N�fT�i��7ui�������F�v��QK���������7�֮�z{�g|+(�8�f=����7�9:)�0!2h�)�o'��BYv��I5���a�������n���v32������¦g�|�Ϫa�-sy5͊��e	�c�*_�Jvq�H���t3n*�:��[QT�h���� �j���*��0j�[��P9�b�V�z5NSa +9KJ�Z��E�Yk�����=���s���Q.����aZ~�r�����-���]w����������顉�qJ�����[a�+�g�$Z��L�Bڇp�C#�7���w�V�@[�8��_+��#��-N���to,qvn�H���T��Ub��X�)�Z���hQ1���5U�^�^���l��N�Ѭ�[�����T��qk��Z%;7�RR�x��OQ縤��b�lH�6|���ߌ����U���/o���?-�Zttl��͛��͙B��2�-���V�?�ĸE]�Eگ7Y���,j�fO���J�M�kC�2�uU錖�"\�j|5��u�K���g����eS.0��	p(�#�FDm�*��wi����������=�4:2J'��ě/�Ї��s���?��/��������hxD�����p�V�^n�x0�N�!�HA�L����l�Mid���;lZ O����uuus�9Ӷh"3Bs��Q&�a���g��3rd�6�?f�B���b�8�ر��n!46Zq�4)����;���*�<Mwv]�^S��n^o�sum�4��C�u�[��k��[�6Z9Ūc)Ɨ� ��~��k?CqnS�\��]��M��3�G/U��*Q��l.KV�xA�c��$l����OdhтE448��wvtr|Z�C��D^�np�̸֤����M��S����qk�wψ���`̅Դx?��Cc�4>6�K/��-7l���t��]�{���|����x�M'��,�Y��K���n��T�[*@/�U�2q�%;;������.Zēi�޽�r,q#�#�����2����� yV�:�
S�D$q�����4�z�:
wl�*INAQ=���<U�E�fs�T�BUl�&�fk�eM�`�њ���ъ�����ܸ�L8y�q����r|i���&c���V���nz���H�I��-=S���U��(2�Vx�,��i�W��]�>P��3���)Ց���Fڠ9=}444D��=40�#�4'ilt����U�R:�	|;S���2��LfhB�3;����Vl�������JnϺ-��8(��'�O���ϱ�&�t�$�8��8w_+@�P�Nf&itl����������l�3��dG}ծ�}xt�z�琝N \�J����"���^@�i�cl���h�Չ��j\���y�����kaKsީDIW�2n��;�zϧ�v�Q�.�j5��u���
�_�Uq�b�RVc7[R�����#��|�Z�T��)Ud��JF���|�=��<�{��``ֿd?E�(��=)��� ��,�;<����o|�a������.���2S��L�)Բ�5A M���蠥K�Ѳ��h�1����-�9��?-&�Yw�[�t��N>pxx�v��C}����e�k��av�gN��Sf��r� t}�Sv�9���J�-�
��R #]U��N,
ƨ�M<%� ,��Z9U�'ٚ�u'����L��7�}b׻�큛f���l�W�W��NZ1~l���8�\��_W��B�qt4��0���
�	3k�[(7��UȠ$C��� >۾���5�l�^�/X��0ǆGhd��c�����֦c�t����Ӫ��hܟl{e���kn���t&���H��[�����={���Ic�WzsP��2j�k[&��o�2��b�S(�kb�T��hq!U�nCWӨh����J<��.��i�*5	Y]UA�7�l:pӫ6�#I)��dT*��IŸ�!m�����&?_�P�h����
�7w2G^�G��s�B���2���mԿ���h!�+���n�a���n~��P�m����'6m����O��~�O=M{�즹s�QgG����>q)"�(+§@yP��4Ot��9AaC��^Q}�ɪR%#�I�x��g�㼩�_�q�U�Yz���i�?��h2M�x��1��G��'�����[�����h�M�~]ƍk��i�U���8!B��p�����4�s����x�������M����9����D�S�vnR�z�	'�������_��/�u�'7-���\F/���F�^�h1��Y�=*:�smx����>��� JU���P���c�#�+����k�N����_�ꈮ�&m4��L�����?��Q�o#�7��6��{�i��F�h���ŐWF�y���`p�w�ذ� ��%�am��A�h��۷����]w޲�+�ziNo?���+p�x����q�'n����:涛6o���_��\:�����W�В�PVt���`�����W1b���T�20Sl���n��v%�i�l�L�R=�fvvj��ꞈ57>��G'M�>X5��M�眢?i�������\U�h��Jjfu��6�l�T*�;�i�`�a�Pf�	q`�/��/����/|��#�z#�ig�&ep�)�_����_������|���Λ�QOoM��a|n��Ϲ��5��7jx��c�J�%������ޗ� �a��ҌӦ�݁������25�2�|b�mGs��e,��)��7����O���86�+[%��{ڪR��G�컃A�Zm��5Q�(�C��tG; �s9����M\����������PE�����>���狟�c�ŗ^:ҿ`	��	��e޼����?|南\t�?t�~���y��͟�K�C#������D� �::;J�}�aH��fL� ͚�຺�҉$�H"�$�l�����l��);9�&E L$�C�\��wR_o/����3����N|ˆM[�<���7�L��q��I�~����?��������#ƁK�9B~���vS_w��-�];_��ή��is��\���'�fK�	#��3� �DI�9���5�̘Z�^�-v	xSxU�Y�l�����*;�#G��� t��n&w�%�����4�f��ٸ��-7ߚ�f��4��rت�;>u��/9y��_�妛���o?�^�˗�si�� ��K�L��k�jюIN��ߍV�6ZU�l�V��X�90�m?��`�yp0Z��=o��?���f{U�pi��Ie#9��)��)7� ,l��tw��9q�F(V�&�40�ݳ�8e�[n}�R�ڙ"3�Iy�i�����G����w_s�����ew#22��j�i<7��R�*�2��1�"v�U)G�F�����V�f8S��rP1�F����K$��mS�ۛ�[b�_�bh�#���ϰWh��C뻼.��f�Y���$�J$K�r�Ḝ�k�\\���=#o�t�×^v���4�eF7�~+Vf����x׻�u�ݟ�����?~���K8��%hK��r�	��zt� ���ȳ����zMfL�^՟H"�T�r��pF ��ׅ���-:9����I�l���$�#�{�Ww�gŊ�������y��h�ȌnRNx۩�V��=����}𪫷��r������C"y���`�$���*K�N(i�*Jy��d�b66�A"�������&�f���9܏a]ߣ����Z���Qޣ��`���r�L�+J�p������y�9�5g�&�5��p���+?����qں��y���zx��D��N#On��^�~L�A�i��\Hf$�-ǃ�>s΢�U�e���kG��� l�x�����a̔�p3Y�d�?�\�	`5�7�_�1A�P�3�H�%�� ��v�A�F[��Ə}��{�����W�:�f��*�&e�CW����G����_��g�>����{߃�t�x��cڿ��Ɔ���Բ,�gs�A��egW';7�����㝦�5#����jU��F�jNAͅ[7����9g���D6x���5+���Q�mv��l	R���y����i���A�_'� p"��ˆ3]t�9߽�K6�Z�꥕���,3{UR���?���\��O<v�����#�ο�o~��Ό���Ҙ��e����R��� v�1���x W�
1�����\w�c��l�|�3ƚ9�[^l]�9�g��Ub+x�ɪ�J������Iw��d���i���~��n����k�^x�E�rʩ�Z��IJ�eV����k�=^����o������s��c��5�޽�v����QJ�Yd��:>6�o:�Iv��k�*��kzw�\���ŏ^��%v�����Se����V�]��=W����PҴ��V|Ą�ɨ����T3�C�F�|��U]��Z����(�}���D�t�_�z�a[n��!X*>E���
`�N�|�R�j`����~�e�����A�*�?"��|ޥ��4�� Z~���|��x�R:�բ�4%R.��%eJ�h�T    IEND�B`�PK   ���XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   ���X�$�  �3     jsons/user_defined.json�Z�n��}A�.�������ڛ¨�	�$(�0ÙaLT&�L�y��L�i/)�N��o��D��s/��;s9����u��̛M�~�!ˋ����Pm�p�G6Mڞ�������˥�m�}�lnҦ������:�-��p���X7��zѡ���O2�ڄ�<��s�E �eH��e�"N�BgJ���Ƹ��ga�|]o3{8�"w𝇠�L{�10ؤ(�<EN:'�!��,Yo�u^�Y9?�4/�۳|�^ُ��
�nN.��p��O/��O,aS�؎DS��H�8�Wu�:Y{B���<�W-&%	��#"����o���)+�z~RW�ʦ�� ��짲��2��C&Eٍ��a��0�f���!���b<
�r@�r�=�W[j�+��g8T��P����;�o�)��޲�v����]5�_]I.�.Ftv��
~����n�ϋ��v}�M��7�&OW��X�5]�CnG`,�-�̺��B�E�?�m�)�Pԛ'� �'we����z�SDS�!n�DF�	��XZ�ӝl�]o�� ҭ}.J��V�+����Yw��}�W���G�8z��+�^��x�3��P���ٕ�E���~��ʣ�E���s�*�"�/CJS�h ,��.L�gh���#�,x�4��3�w�2������%!C�Ad±��pӀ�L4WD-�I���M{ƛ���B���(�#}����(�F��C���C9�޷��_��9ۇ��˳(S�J:Nk'�m=� C�E6(	+pㅒ;nLi`P6}a\��̀�!�U���9=}$��M�GƦ�[Pqj�D�BIe�2���B��i�b����Im%
^p��4 �!(hǝ�R����~Ȃ�J�����MY�z�w�S���Gٔ�I��x�B�ž�Ds�(`�Zh�	���j�:�8@m��C�a���� �����g���Y���OZ|.���튋�ǋ<���]���GW1�8���sO0�S��c0$Lpwa3���lf�3I�������P��<�2�pW��r7_�x/7������'�`A�~

?v"@(�\LSR!��HE>.��J���T�r�Qz2'81�@=����w*���|o�9��<�h�'��=�%)�A8dS(�2�*{W߿avH�D�����fU�׳��7�5ቦ�O0�[V�ɋr����#������GSW�j�3�0��C-�P�L����0m��#
&��Ɩ��S���b�A��� �+dp@Xg�JY�.m��N���)�}+F��!�Rrx"L��g������_��?��>R���<;���2lB}��NF��r��(*(T1�)��:
���#��j�T���8
���(�%�4}�<Ɯ(a�8�/�8�@�%��K6:�\�������R⨿�}=��cA��e&'���d2�)��2@җ�q�Sb%}a{F&���ᱰ�B�EK���-;�/t�h�HX3�:P�t$�G�k�s�T5���%��r�/��Ġ���[,u��@�⑨���KD�����.�:..6P�T$*[�?���d�kF��m����L�0wO3j��e߱�Z��@)�'��B��fq3�|S��{�?�<��9u�F��2�yPH+P��\9턍];Y�,w#�S	h�P*�@�P̌�t�n�h��j;�]�a!&����Ӟ����L� �α�ǰ�|ٴ���|�[��@r0�{z��ߏ�����]����x�������/��!_~(�*a��uܹ����ڤ�8��!���ݷ�3m��~�?�D����\6�i�fϳ�϶𛇜ė	�XȨX_�7`��¡uC���{h˘ XQn�~�jGG8:����pt��#��C���&T�v5{�n��m�y��݉����� ��vcLȐ�Z�`u�Y���Xr��6㰌HiҾ�pq�6>CY걂CXZ��r�8�hʐ!�'#p���4�$X���H~����|�-���T����z$#	&\��J%���jڔ&����D����L`�:и�G���0�V�>Hћ>_�PK
   ���X�v�[E7  `�                  cirkitFile.jsonPK
   ���X��g  n  /             r7  images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.pngPK
   ���X�j�� 7q /             &P  images/3afa6c98-60d7-4a37-9aec-be07fd386e0e.pngPK
   ���XhT���� ċ /             �5 images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.pngPK
   C��X�y�H$  �G  /             `� images/81d9366d-a3a2-4692-b3d3-374cda370674.pngPK
   ���Xd��  �   /             �	 images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   ��Xք|� t� /             '	 images/83f16691-8d82-4f83-89df-fbd07d8206a1.pngPK
   ���X	�\  \  /             ��
 images/898ac7d1-13d0-4a1b-8b5c-ab7066f4327a.pngPK
   C��X o
7  �%  /             } images/8bec88c5-4482-4569-926a-ae76def9d576.pngPK
   ���X	��#u } /             # images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   C��X����?  [G  /             q� images/b3b368a6-ed54-49be-b991-e8c4c6667997.pngPK
   ���X$7h�!  �!  /             l� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   C��X��iP  K  /             �� images/e6075517-c690-4ca2-aabd-cadc5d2d7233.pngPK
   ��X�3S�u� �� /             L images/ec43f2b3-9126-4f13-83de-62ba1ea97088.pngPK
   ���XP��/�  ǽ  /             � images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   ���X�$�  �3               `h jsons/user_defined.jsonPK      �  �p   